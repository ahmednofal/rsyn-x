module cpu ( gnd, vdd, clk, reset, DI_0_, DI_1_, DI_2_, DI_3_, DI_4_, DI_5_, DI_6_, DI_7_, IRQ, NMI, RDY, AB_0_, AB_1_, AB_2_, AB_3_, AB_4_, AB_5_, AB_6_, AB_7_, AB_8_, AB_9_, AB_10_, AB_11_, AB_12_, AB_13_, AB_14_, AB_15_, DO_0_, DO_1_, DO_2_, DO_3_, DO_4_, DO_5_, DO_6_, DO_7_, WE);

input gnd, vdd;
input clk;
input reset;
input DI_0_;
input DI_1_;
input DI_2_;
input DI_3_;
input DI_4_;
input DI_5_;
input DI_6_;
input DI_7_;
input IRQ;
input NMI;
input RDY;
output AB_0_;
output AB_1_;
output AB_2_;
output AB_3_;
output AB_4_;
output AB_5_;
output AB_6_;
output AB_7_;
output AB_8_;
output AB_9_;
output AB_10_;
output AB_11_;
output AB_12_;
output AB_13_;
output AB_14_;
output AB_15_;
output DO_0_;
output DO_1_;
output DO_2_;
output DO_3_;
output DO_4_;
output DO_5_;
output DO_6_;
output DO_7_;
output WE;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf5) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf4) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf3) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf2) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf1) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf0) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_980_), .Y(_980__bF_buf4) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_980_), .Y(_980__bF_buf3) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(_980_), .Y(_980__bF_buf2) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_980_), .Y(_980__bF_buf1) );
	BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_980_), .Y(_980__bF_buf0) );
	BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .Y(_1100__bF_buf3) );
	BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .Y(_1100__bF_buf2) );
	BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .Y(_1100__bF_buf1) );
	BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .Y(_1100__bF_buf0) );
	BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_929_), .Y(_929__bF_buf4) );
	BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_929_), .Y(_929__bF_buf3) );
	BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_929_), .Y(_929__bF_buf2) );
	BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_929_), .Y(_929__bF_buf1) );
	BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_929_), .Y(_929__bF_buf0) );
	BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf7) );
	BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf6) );
	BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf5) );
	BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf4) );
	BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf3) );
	BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf2) );
	BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf1) );
	BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf0) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .Y(_1789__bF_buf3) );
	BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .Y(_1789__bF_buf2) );
	BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .Y(_1789__bF_buf1) );
	BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .Y(_1789__bF_buf0) );
	BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_928__bF_buf4) );
	BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_928__bF_buf3) );
	BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_928__bF_buf2) );
	BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_928__bF_buf1) );
	BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_928__bF_buf0) );
	BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_953_), .Y(_953__bF_buf4) );
	BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_953_), .Y(_953__bF_buf3) );
	BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_953_), .Y(_953__bF_buf2) );
	BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_953_), .Y(_953__bF_buf1) );
	BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_953_), .Y(_953__bF_buf0) );
	BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_578__bF_buf4) );
	BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_578__bF_buf3) );
	BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_578__bF_buf2) );
	BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_578__bF_buf1) );
	BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_578__bF_buf0) );
	BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf8) );
	BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf7) );
	BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf6) );
	BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf5) );
	BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf4) );
	BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf3) );
	BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf2) );
	BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf1) );
	BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf0) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_939_), .Y(_939__bF_buf3) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_939_), .Y(_939__bF_buf2) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_939_), .Y(_939__bF_buf1) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_939_), .Y(_939__bF_buf0) );
	BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .Y(_1077__bF_buf3) );
	BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .Y(_1077__bF_buf2) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .Y(_1077__bF_buf1) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .Y(_1077__bF_buf0) );
	BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .Y(_1065__bF_buf3) );
	BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .Y(_1065__bF_buf2) );
	BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .Y(_1065__bF_buf1) );
	BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .Y(_1065__bF_buf0) );
	BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf4) );
	BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf3) );
	BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf2) );
	BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf1) );
	BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf0) );
	BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf4) );
	BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf3) );
	BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf2) );
	BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf1) );
	BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf0) );
	BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1509__bF_buf4) );
	BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1509__bF_buf3) );
	BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1509__bF_buf2) );
	BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1509__bF_buf1) );
	BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1509__bF_buf0) );
	BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(_979_), .Y(_979__bF_buf3) );
	BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(_979_), .Y(_979__bF_buf2) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_979_), .Y(_979__bF_buf1) );
	BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(_979_), .Y(_979__bF_buf0) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .Y(_924_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(state_4_), .Y(_925_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_926_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_927_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf5), .B(_926_), .C(_927_), .Y(_928_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_928__bF_buf4), .Y(_929_) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .Y(_930_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_4_), .Y(_932_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(DI_4_), .Y(_933_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_932_), .C(_933_), .Y(DIMUX_4_) );
	INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_4_), .Y(_934_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(I), .Y(_935_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(IRQ), .Y(_936_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(NMI_edge), .Y(_937_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_937_), .Y(_938_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(NMI_edge), .C(_938_), .Y(_939_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(IRHOLD_4_), .C(_939__bF_buf3), .Y(_940_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_934_), .C(_940_), .Y(_941_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_3_), .Y(_942_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_3_), .Y(_943_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(DI_3_), .Y(_944_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_943_), .C(_944_), .Y(DIMUX_3_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(DIMUX_3_), .Y(_945_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_942_), .C(_945_), .Y(_946_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_939__bF_buf2), .B(_946_), .Y(_947_) );
	MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(DI_2_), .B(DIHOLD_2_), .S(RDY_bF_buf3), .Y(_948_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_2_), .Y(_949_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_948_), .C(_949_), .Y(_950_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_939__bF_buf1), .Y(_951_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_947_), .Y(_952_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(I), .B(_936_), .C(_937_), .Y(_953_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_1_), .Y(_954_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(DI_1_), .Y(_955_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_954_), .C(_955_), .Y(DIMUX_1_) );
	MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .B(IRHOLD_1_), .S(_930_), .Y(_956_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_953__bF_buf4), .Y(_957_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_0_), .Y(_958_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(DI_0_), .Y(_959_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_958_), .C(_959_), .Y(DIMUX_0_) );
	MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(IRHOLD_0_), .S(_930_), .Y(_960_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf3), .B(_960_), .Y(_961_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_961_), .Y(_962_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_962_), .Y(_963_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_946_), .C(_939__bF_buf0), .Y(_964_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_4_), .Y(_965_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_965_), .C(_953__bF_buf2), .Y(_966_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(DIMUX_4_), .C(_966_), .Y(_967_) );
	MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(DI_7_), .B(DIHOLD_7_), .S(RDY_bF_buf7), .Y(_968_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_7_), .Y(_969_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_968_), .C(_969_), .Y(_970_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_939__bF_buf3), .Y(_971_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_971_), .Y(_972_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_972_), .Y(_973_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_973_), .Y(_974_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_963_), .C(_974_), .Y(_975_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_976_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_976_), .Y(_977_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_978_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_977_), .Y(_979_) );
	INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf4), .Y(_980_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(_981_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_981_), .Y(_982_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_983_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_982_), .Y(_984_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf3), .B(_984_), .Y(_985_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf3), .B(_980__bF_buf4), .C(_985_), .Y(_986_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(state_4_), .Y(_987_) );
	INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_987_), .Y(_988_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .Y(_989_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_989_), .Y(_990_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_991_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_992_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_992_), .Y(_993_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_993_), .Y(_994_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_979__bF_buf2), .C(_994_), .Y(_995_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_986_), .Y(_996_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf1), .Y(_997_) );
	INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(_998_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_998_), .Y(_999_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_998_), .Y(_1000_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(state_1_), .C(_927_), .Y(_1001_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001_), .Y(_1002_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_999_), .C(_1002_), .Y(_1003_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_976_), .C(_991_), .Y(_1004_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_989_), .Y(_1005_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1005__bF_buf4), .Y(_1006_) );
	INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_1007_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_1007_), .Y(_1008_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_1008_), .Y(_1009_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1009_), .Y(_1010_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1006_), .C(_1010_), .Y(_1011_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_1011_), .Y(_1012_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_996_), .C(_1012_), .Y(_1013_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_977_), .Y(_1014_) );
	NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .C(_991_), .Y(_1015_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1015_), .Y(_1016_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1014_), .C(_1016_), .Y(_1017_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_990_), .Y(_1018_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_984_), .Y(_1019_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf3), .B(_1014_), .Y(_1020_) );
	INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .Y(_1021_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(store), .Y(_1022_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1022_), .Y(_1023_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1023_), .C(RDY_bF_buf2), .D(_1021_), .Y(_1024_) );
	AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_1025_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_1025_), .Y(_1026_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .Y(_1027_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf2), .B(_1027_), .Y(_1028_) );
	INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(write_back), .Y(_1029_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(RDY_bF_buf1), .C(_1022_), .Y(_1030_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1028_), .Y(_1031_) );
	NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1018_), .C(_1024_), .Y(_1032_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_995_), .Y(_1033_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(RDY_bF_buf0), .C(_1033_), .Y(_1034_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_1034_), .C(_1032_), .Y(_1035_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_929__bF_buf4), .C(_1035_), .Y(_1036_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf1), .B(_956_), .Y(_1037_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_961_), .Y(_1038_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_1038_), .Y(_1039_) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(DIMUX_4_), .Y(_1040_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_965_), .C(_1040_), .Y(_1041_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_1041_), .C(_939__bF_buf2), .Y(_1042_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_5_), .Y(_1043_) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(DI_5_), .Y(_1044_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1043_), .C(_1044_), .Y(DIMUX_5_) );
	MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .B(IRHOLD_5_), .S(_930_), .Y(_1045_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf0), .B(_1045_), .Y(_1046_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_6_), .Y(_1047_) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(DI_6_), .Y(_1048_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1047_), .C(_1048_), .Y(DIMUX_6_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_6_), .Y(_1049_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_1049_), .C(_953__bF_buf4), .Y(_1050_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(DIMUX_6_), .C(_1050_), .Y(_1051_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1046_), .Y(_1052_) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1052_), .Y(_1053_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1039_), .Y(_1054_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_990_), .C(_1008_), .Y(_1055_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .Y(_1056_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf6), .B(_1056_), .C(_929__bF_buf3), .D(_1054_), .Y(_1057_) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1010_), .Y(_1058_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(store), .C(RDY_bF_buf4), .Y(_1059_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1059_), .C(_1058_), .Y(_1060_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .Y(_1061_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1061_), .C(_1036_), .Y(_1062_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_994_), .Y(_1063_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_946_), .C(_939__bF_buf1), .Y(_1064_) );
	INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf2), .Y(_1065_) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_939__bF_buf0), .B(_950_), .Y(_1066_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1065__bF_buf3), .Y(_1067_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_1063_), .C(_1064_), .D(_1067_), .Y(_1068_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf2), .B(_1001_), .C(RDY_bF_buf3), .Y(_1069_) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_1025_), .Y(_1070_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf1), .B(_1070_), .Y(_1071_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_1071_), .C(_1069_), .Y(_1072_) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1068_), .Y(_1073_) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1008_), .Y(_1074_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1074_), .Y(_1075_) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_976_), .Y(_1076_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_1076_), .Y(_1077_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_1077__bF_buf3), .Y(_1078_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1078_), .C(RDY_bF_buf1), .Y(_1079_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1075_), .C(_1079_), .Y(_1080_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1074_), .Y(_1081_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1078_), .C(RDY_bF_buf8), .Y(_1082_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1081_), .C(_1082_), .Y(_1083_) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1083_), .Y(_1084_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1073_), .Y(_1085_) );
	NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_981_), .C(_992_), .Y(_1086_) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_1086_), .Y(_1087_) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_1007_), .Y(_1088_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1088_), .Y(_1089_) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_1089_), .Y(_1090_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .Y(_1091_) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1091_), .Y(_1092_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1087_), .C(_1092_), .Y(_1093_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(state_3_), .C(_1025_), .Y(_1094_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf0), .B(_1094_), .Y(_1095_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .Y(_1096_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_1097_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_1097_), .Y(_1098_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_981_), .Y(_1099_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf1), .B(_1098_), .C(_1099_), .Y(_1100_) );
	MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1100__bF_buf3), .S(_924__bF_buf3), .Y(_1101_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(_1093_), .Y(_1102_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1094_), .C(_924__bF_buf2), .Y(_1103_) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1099_), .Y(_1104_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf4), .B(_1104_), .Y(_1105_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_1105_), .C(_1103_), .Y(_1106_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf0), .B(_1008_), .C(_1098_), .Y(_1107_) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(backwards), .Y(_1108_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .Y(_1109_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_1109_), .C(RDY_bF_buf4), .Y(_1110_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf4), .B(_1074_), .Y(_1111_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1111_), .C(_1110_), .Y(_1112_) );
	AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1106_), .Y(_1113_) );
	AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1113_), .Y(_1114_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_924__bF_buf0), .Y(_1115_) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1026_), .Y(_1116_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_1116_), .C(_1115_), .D(_1033_), .Y(_1117_) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1026_), .Y(_1118_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(state_1_), .C(_978_), .Y(_1119_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1119_), .C(RDY_bF_buf2), .Y(_1120_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1118_), .C(_1120_), .Y(_1121_) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1117_), .Y(_1122_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_999_), .C(_1098_), .Y(_1123_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .Y(_1124_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1070_), .C(_924__bF_buf6), .Y(_1125_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1124_), .C(_1125_), .Y(_1126_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf3), .B(_1026_), .C(_924__bF_buf4), .Y(_1127_) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf2), .B(_1119_), .Y(_1128_) );
	OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1128_), .C(_1127_), .Y(_1129_) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1126_), .Y(_1130_) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1122_), .Y(_1131_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1114_), .C(_1131_), .Y(_1132_) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_979__bF_buf0), .Y(_1133_) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_1133_), .Y(_1134_) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_939__bF_buf3), .B(_970_), .Y(_1135_) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_967_), .Y(_1136_) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1136_), .Y(_1137_) );
	INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_3_), .Y(_1138_) );
	OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(IRHOLD_3_), .C(_939__bF_buf2), .Y(_1139_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_1138_), .C(_1139_), .Y(_1140_) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1140_), .Y(_1141_) );
	OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf3), .B(_960_), .C(_957_), .Y(_1142_) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1142_), .Y(_1143_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf1), .B(_1137_), .C(_1143_), .Y(_1144_) );
	AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1134_), .Y(_1145_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf5), .B(_977_), .C(_1008_), .Y(_1146_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .Y(_1147_) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1039_), .Y(_1148_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_1147_), .C(_929__bF_buf0), .D(_1148_), .Y(_1149_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_926_), .C(_987_), .Y(_1150_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .Y(_1151_) );
	OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_979__bF_buf3), .C(_924__bF_buf0), .Y(_1152_) );
	OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_1151_), .C(_1152_), .Y(_1153_) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_926_), .Y(_1154_) );
	NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1154_), .Y(_1155_) );
	OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf4), .B(_979__bF_buf2), .C(_924__bF_buf6), .Y(_1156_) );
	OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1155_), .C(_1156_), .Y(_1157_) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1153_), .Y(_1158_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .Y(_1159_) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_1099_), .Y(_1160_) );
	OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1160_), .C(_924__bF_buf4), .Y(_1161_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(state_3_), .C(_926_), .Y(_1162_) );
	NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1162_), .Y(_1163_) );
	OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1163_), .C(_1161_), .Y(_1164_) );
	NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf1), .B(_1160_), .Y(_1165_) );
	NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1165_), .Y(_1166_) );
	NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_1088_), .Y(_1167_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_925__bF_buf4), .C(_924__bF_buf2), .Y(_1168_) );
	OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1166_), .C(_1164_), .Y(_1169_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_925__bF_buf3), .C(_926_), .Y(_1170_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .Y(_1171_) );
	OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf0), .B(_979__bF_buf1), .C(_924__bF_buf1), .Y(_1172_) );
	OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_1171_), .C(_1172_), .Y(_1173_) );
	OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1160_), .C(_924__bF_buf7), .Y(_1174_) );
	NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1162_), .Y(_1175_) );
	OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf6), .B(_1175_), .C(_1174_), .Y(_1176_) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1017_), .Y(_1177_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1176_), .C(_1177_), .Y(_1178_) );
	NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1169_), .Y(_1179_) );
	AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1159_), .Y(_1180_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_1180_), .C(_1145_), .Y(_1181_) );
	NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1132_), .C(_1062_), .Y(_1182_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .Y(_919_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .Y(_1183_) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1046_), .Y(_1184_) );
	NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1184_), .Y(_1185_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf4), .B(_1185_), .C(_1143_), .Y(_1186_) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1124_), .Y(_1187_) );
	OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1001_), .C(_924__bF_buf4), .Y(_1188_) );
	OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1116_), .C(_1188_), .Y(_1189_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1189_), .C(_1186_), .Y(_1190_) );
	NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_961_), .Y(_1191_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_957_), .C(_1191_), .Y(_1192_) );
	NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1192_), .Y(_1193_) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1077__bF_buf2), .Y(_1194_) );
	NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1160_), .Y(_1195_) );
	OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1195_), .C(RDY_bF_buf8), .Y(_1196_) );
	OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1194_), .C(_1196_), .Y(_1197_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(_929__bF_buf3), .C(_1197_), .Y(_1198_) );
	NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf4), .B(_1001_), .Y(_1199_) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_1199_), .Y(_1200_) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_962_), .Y(_1201_) );
	NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1201_), .Y(_1202_) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf2), .B(_1202_), .Y(_1203_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1203_), .C(_1198_), .Y(_1204_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_953__bF_buf2), .Y(_1205_) );
	NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1205_), .Y(_1206_) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1051_), .Y(_1207_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1208_) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1206_), .Y(_1209_) );
	NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1209_), .Y(_1210_) );
	AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_1105_), .C(_929__bF_buf1), .D(_1210_), .Y(_1211_) );
	NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_971_), .Y(_1212_) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1206_), .Y(_1213_) );
	NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1213_), .Y(_1214_) );
	AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_1091_), .C(_929__bF_buf0), .D(_1214_), .Y(_1215_) );
	NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_1146_), .Y(_1216_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(Z), .Y(_1217_) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_1217_), .Y(_1218_) );
	OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(C), .C(_1218_), .Y(_1219_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(V), .Y(_1220_) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_1220_), .Y(_1221_) );
	OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(N), .B(cond_code_1_), .C(_1221_), .Y(_1222_) );
	MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(_1222_), .S(cond_code_2_), .Y(_1223_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(cond_code_0_), .Y(_1224_) );
	OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1078_), .C(_924__bF_buf6), .Y(_1225_) );
	OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1056_), .C(_1225_), .Y(_1226_) );
	OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1107_), .C(_1226_), .Y(_1227_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1216_), .C(_1227_), .Y(_1228_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1211_), .C(_1215_), .Y(_1229_) );
	NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1204_), .C(_1229_), .Y(_1230_) );
	NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1119_), .Y(_1231_) );
	NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1201_), .Y(_1232_) );
	AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_1231_), .C(_929__bF_buf4), .D(_1232_), .Y(_1233_) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_1097_), .Y(_1234_) );
	NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1088_), .Y(_1235_) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf2), .B(_1235_), .Y(_1236_) );
	INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf2), .Y(_1237_) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1237_), .Y(_1238_) );
	OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_1236_), .C(_1238_), .Y(_1239_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .Y(_1240_) );
	NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1119_), .Y(_1241_) );
	OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_979__bF_buf0), .C(RDY_bF_buf5), .Y(_1242_) );
	OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1241_), .C(_1242_), .Y(_1243_) );
	OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1240_), .C(_1243_), .Y(_1244_) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1239_), .Y(_1245_) );
	OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf1), .B(_956_), .C(_961_), .Y(_1246_) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_1140_), .Y(_1247_) );
	OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1141_), .C(_1247_), .Y(_1248_) );
	NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1065__bF_buf2), .Y(_1249_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1249_), .C(_1245_), .Y(_1250_) );
	AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1250_), .Y(_1251_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1251_), .C(_1230_), .Y(_920_) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_1008_), .Y(_1252_) );
	OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf4), .B(_1252_), .C(_924__bF_buf1), .Y(_1253_) );
	OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_1118_), .C(_1253_), .Y(_1254_) );
	NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_1033_), .Y(_1255_) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_1256_) );
	NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1076_), .Y(_1258_) );
	OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_1235_), .C(_990_), .Y(_1259_) );
	OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_1074_), .C(_1259_), .Y(_1260_) );
	NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1154_), .Y(_1261_) );
	NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1252_), .Y(_1262_) );
	NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1262_), .Y(_1263_) );
	OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf3), .B(_1014_), .C(_1263_), .Y(_1264_) );
	OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1264_), .C(_1255_), .Y(_1265_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1266_) );
	INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .Y(_1267_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_1109_), .C(_1267_), .Y(_1268_) );
	OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_928__bF_buf3), .C(_1268_), .Y(_1269_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1216_), .C(_1269_), .Y(_1270_) );
	AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1270_), .Y(_1271_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_967_), .C(_1039_), .Y(_1272_) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1143_), .Y(_1273_) );
	OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1201_), .C(_1273_), .Y(_1274_) );
	NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1274_), .Y(_1275_) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1143_), .Y(_1276_) );
	OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1213_), .C(_1276_), .Y(_1277_) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_947_), .Y(_1278_) );
	NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1278_), .Y(_1279_) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1279_), .Y(_1280_) );
	OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1213_), .C(_1280_), .Y(_1281_) );
	NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1281_), .B(_1277_), .Y(_1282_) );
	NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1141_), .Y(_1283_) );
	AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_973_), .C(_967_), .D(_1283_), .Y(_1284_) );
	OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1140_), .C(_929__bF_buf3), .Y(_1285_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .Y(_1286_) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1284_), .Y(_1287_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1248_), .C(_1287_), .Y(_1288_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1282_), .C(_1288_), .Y(_1289_) );
	NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1142_), .Y(_1290_) );
	OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1184_), .C(_972_), .Y(_1291_) );
	OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf0), .B(_960_), .C(_1037_), .Y(_1292_) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1292_), .Y(_1293_) );
	NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1247_), .Y(_1294_) );
	AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1293_), .Y(_1295_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1291_), .C(_1295_), .Y(_1296_) );
	NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1141_), .Y(_1297_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1136_), .C(_1297_), .Y(_1298_) );
	OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf4), .B(_1045_), .C(_967_), .Y(_1299_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .Y(_1300_) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1300_), .Y(_1301_) );
	NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1301_), .Y(_1302_) );
	INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_6_), .Y(_1303_) );
	OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(IRHOLD_6_), .C(_939__bF_buf1), .Y(_1304_) );
	AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_1303_), .C(_1304_), .Y(_1305_) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1305_), .Y(_1306_) );
	NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1306_), .Y(_1307_) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1290_), .Y(_1308_) );
	OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1209_), .C(_1308_), .Y(_1309_) );
	NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1309_), .Y(_1310_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1298_), .C(_1310_), .Y(_1311_) );
	OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1289_), .C(_1271_), .Y(_1312_) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_927_), .Y(_1313_) );
	NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1313_), .Y(_1314_) );
	OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1094_), .C(RDY_bF_buf0), .Y(_1315_) );
	OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1314_), .C(_1315_), .Y(_1316_) );
	NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1313_), .Y(_1317_) );
	OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1094_), .C(RDY_bF_buf7), .Y(_1318_) );
	OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1317_), .C(_1318_), .Y(_1319_) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .B(_1316_), .Y(_1320_) );
	NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1312_), .Y(_1321_) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1190_), .Y(_1322_) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf6), .B(_1262_), .Y(_1323_) );
	OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf1), .B(_1298_), .C(_1323_), .Y(_1324_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_985_), .Y(_1325_) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(write_back), .B(RDY_bF_buf5), .Y(_1326_) );
	AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1326_), .C(_1028_), .Y(_1327_) );
	AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_924__bF_buf5), .C(_1327_), .Y(_1328_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .Y(_1329_) );
	NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1324_), .Y(_1330_) );
	AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1177_), .Y(_1331_) );
	AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_1126_), .Y(_1332_) );
	AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1228_), .Y(_1333_) );
	AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1149_), .Y(_1334_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1334_), .C(_1330_), .Y(_1335_) );
	NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1322_), .C(_1335_), .Y(_1336_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1336_), .C(_1321_), .Y(_921_) );
	AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1185_), .C(_941_), .D(_1248_), .Y(_1337_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1298_), .C(_1337_), .Y(_1338_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .Y(_1339_) );
	NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1142_), .Y(_1340_) );
	NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1306_), .Y(_1341_) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1340_), .Y(_1342_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1308_), .C(_1342_), .Y(_1343_) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1344_) );
	AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1137_), .C(_1285_), .Y(_1345_) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1344_), .Y(_1346_) );
	NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_1343_), .C(_1346_), .Y(_1347_) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1290_), .Y(_1348_) );
	NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1232_), .Y(_1349_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1296_), .C(_1349_), .Y(_1350_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .Y(_1351_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1347_), .C(_1351_), .Y(_1352_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .Y(_1353_) );
	NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1353_), .Y(_1354_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1271_), .B(_1354_), .C(_1352_), .Y(_1355_) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_952_), .Y(_1356_) );
	NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1356_), .Y(_1357_) );
	OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .B(_1357_), .C(_929__bF_buf2), .Y(_1358_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1328_), .C(_1358_), .Y(_1359_) );
	NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1140_), .Y(_1360_) );
	AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_1151_), .C(_1249_), .D(_1360_), .Y(_1361_) );
	OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf2), .B(_1070_), .C(RDY_bF_buf4), .Y(_1362_) );
	OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1155_), .C(_1362_), .Y(_1363_) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1361_), .Y(_1364_) );
	OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1070_), .C(RDY_bF_buf2), .Y(_1365_) );
	OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1261_), .C(_1365_), .Y(_1366_) );
	OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1170_), .C(_1366_), .Y(_1367_) );
	NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1364_), .Y(_1368_) );
	NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1368_), .C(_1233_), .Y(_1369_) );
	NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf1), .B(_1341_), .C(_1290_), .Y(_1370_) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1175_), .Y(_1372_) );
	AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1372_), .Y(_1373_) );
	OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1074_), .C(RDY_bF_buf8), .Y(_1374_) );
	OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1163_), .C(_1374_), .Y(_1375_) );
	AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1291_), .Y(_1376_) );
	OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1376_), .C(_929__bF_buf0), .Y(_1377_) );
	NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1375_), .C(_1377_), .Y(_1378_) );
	NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1359_), .B(_1369_), .C(_1378_), .Y(_1379_) );
	NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1379_), .C(_1182_), .Y(_1380_) );
	OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf0), .B(_1280_), .C(_1200_), .Y(_1381_) );
	NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_1320_), .C(_1169_), .Y(_1382_) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1126_), .B(_1106_), .Y(_1383_) );
	NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1177_), .Y(_1384_) );
	NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1383_), .Y(_1385_) );
	NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1385_), .C(_1382_), .Y(_1386_) );
	NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1386_), .C(_1381_), .Y(_1387_) );
	NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1215_), .Y(_1389_) );
	NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1389_), .Y(_1390_) );
	NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf3), .B(_1284_), .Y(_1391_) );
	NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1375_), .C(_1370_), .Y(_1392_) );
	NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1392_), .C(_1391_), .Y(_1393_) );
	NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1393_), .C(_1390_), .Y(_1394_) );
	NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_1312_), .Y(_1396_) );
	OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1380_), .C(_1396_), .Y(_922_) );
	NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .B(_1254_), .C(_1061_), .Y(_1397_) );
	NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1080_), .Y(_1398_) );
	NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1397_), .Y(_1399_) );
	NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1385_), .C(_1399_), .Y(_1400_) );
	NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1400_), .Y(_1401_) );
	NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1373_), .C(_1401_), .Y(_1403_) );
	AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1187_), .Y(_1404_) );
	NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1404_), .C(_1211_), .Y(_1405_) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1405_), .Y(_923_) );
	NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1145_), .C(_1215_), .Y(_1407_) );
	AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1243_), .Y(_1408_) );
	NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1408_), .C(_1117_), .Y(_1409_) );
	NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1093_), .Y(_1410_) );
	NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1164_), .C(_1410_), .Y(_1411_) );
	AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(_1316_), .Y(_1412_) );
	NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1366_), .C(_1412_), .Y(_1413_) );
	OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1413_), .Y(_1414_) );
	NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1414_), .Y(_1415_) );
	NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1361_), .C(_1415_), .Y(_1416_) );
	NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1416_), .Y(_1417_) );
	NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1323_), .C(_1417_), .Y(_931_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(C), .Y(_1419_) );
	INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(shift), .Y(_1420_) );
	OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_984_), .B(_1027_), .C(_990_), .Y(_1421_) );
	OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf1), .B(_1014_), .C(_1421_), .Y(_1422_) );
	NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(load_only), .B(_1021_), .Y(_1423_) );
	AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(rotate), .B(_1422_), .C(_1420_), .D(_1423_), .Y(_1425_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(rotate), .Y(_1426_) );
	INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(compare), .Y(_1427_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .Y(_1428_) );
	NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(inc), .C(_1428_), .Y(_1429_) );
	OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1021_), .C(_1429_), .Y(_1430_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1431_) );
	OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf0), .B(_1026_), .C(_1107_), .Y(_1433_) );
	OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1431_), .C(ALU_CO), .Y(_1434_) );
	INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .Y(_1435_) );
	OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf4), .B(_1070_), .C(_1435_), .Y(_1436_) );
	OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1119_), .C(_1087_), .Y(_1437_) );
	NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1437_), .B(_1436_), .Y(_1438_) );
	AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_1077__bF_buf1), .C(_1124_), .Y(_1439_) );
	OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1104_), .C(_1055_), .Y(_1440_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .Y(_1441_) );
	AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1441_), .Y(_1442_) );
	NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1438_), .C(_1442_), .Y(_1443_) );
	AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1430_), .C(_1443_), .Y(_1444_) );
	OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_1425_), .C(_1444_), .Y(ALU_CI) );
	INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(PC_0_), .Y(_1445_) );
	INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .Y(_1446_) );
	NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_1165_), .Y(_1447_) );
	NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1105_), .Y(_1448_) );
	AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1015_), .C(_990_), .D(_1258_), .Y(_1449_) );
	NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_1104_), .Y(_1450_) );
	NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf1), .B(_926_), .C(_1099_), .Y(_1451_) );
	OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1252_), .C(_1451_), .Y(_1452_) );
	NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1452_), .Y(_1453_) );
	NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1448_), .C(_1453_), .Y(_1454_) );
	AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_1086_), .C(_1436_), .Y(_1455_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1456_) );
	AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_1456_), .C(_1133_), .Y(_1457_) );
	NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1457_), .C(_1455_), .Y(_1458_) );
	NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1458_), .Y(_1459_) );
	NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1459_), .Y(_1460_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_1146_), .C(_1446_), .D(_1460_), .Y(ALU_BI_0_) );
	INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(PC_1_), .Y(_1461_) );
	INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .Y(_1462_) );
	OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1146_), .C(_1462_), .D(_1460_), .Y(ALU_BI_1_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(DIMUX_2_) );
	INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .Y(_1463_) );
	OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1146_), .C(_948_), .D(_1460_), .Y(ALU_BI_2_) );
	INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .Y(_1464_) );
	OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1146_), .C(_1138_), .D(_1460_), .Y(ALU_BI_3_) );
	INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .Y(_1465_) );
	OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_1146_), .C(_934_), .D(_1460_), .Y(ALU_BI_4_) );
	INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .Y(_1466_) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .Y(_1467_) );
	OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1146_), .C(_1467_), .D(_1460_), .Y(ALU_BI_5_) );
	INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .Y(_1468_) );
	OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1146_), .C(_1303_), .D(_1460_), .Y(ALU_BI_6_) );
	INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_968_), .Y(DIMUX_7_) );
	INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .Y(_1469_) );
	OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1146_), .C(_968_), .D(_1460_), .Y(ALU_BI_7_) );
	NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_1077__bF_buf0), .Y(_1470_) );
	NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf1), .B(_1470_), .C(_1236_), .Y(_1471_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .Y(_1472_) );
	NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .B(_1455_), .Y(_1473_) );
	OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1026_), .C(_1146_), .Y(_1474_) );
	INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .Y(_1475_) );
	NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(ABH_0_), .B(_925__bF_buf0), .C(_1077__bF_buf3), .Y(_1476_) );
	OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1475_), .C(_1476_), .Y(_1477_) );
	AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_0_), .C(_1477_), .Y(_1478_) );
	INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf2), .Y(_1479_) );
	OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1005__bF_buf4), .C(_980__bF_buf3), .D(_1001_), .Y(_1480_) );
	OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf2), .B(_1119_), .C(_1150_), .Y(_1481_) );
	OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1481_), .Y(_1482_) );
	AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_1_), .B(_1479_), .C(_1482_), .Y(_1483_) );
	OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1313_), .C(_1000__bF_buf4), .D(_1119_), .Y(_1484_) );
	AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_1313_), .C(_1000__bF_buf3), .Y(_1485_) );
	NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_1485_), .Y(_1486_) );
	OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1005__bF_buf2), .C(_980__bF_buf1), .D(_1094_), .Y(_1487_) );
	AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_1089_), .C(_1487_), .Y(_1488_) );
	NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1123_), .C(_1055_), .Y(_1489_) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .Y(_1490_) );
	NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1486_), .C(_1490_), .Y(_1491_) );
	OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf0), .B(_1313_), .C(src_reg_1_), .Y(_1492_) );
	OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1491_), .C(_1483_), .Y(_1493_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__0_), .Y(_1494_) );
	AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_925__bF_buf5), .C(_999_), .D(_1089_), .Y(_1495_) );
	NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_1097_), .C(_991_), .Y(_1496_) );
	AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1496_), .C(_990_), .D(_1089_), .Y(_1497_) );
	NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1497_), .C(_1495_), .Y(_1498_) );
	AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_999_), .C(_925__bF_buf4), .D(_1086_), .Y(_1499_) );
	OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1167_), .C(_990_), .Y(_1500_) );
	NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .B(_1449_), .C(_1500_), .Y(_1501_) );
	NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1498_), .Y(_1502_) );
	OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf4), .B(_1313_), .C(src_reg_0_), .Y(_1503_) );
	NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(_1481_), .C(_1480_), .Y(_1504_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .Y(_1505_) );
	NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_0_), .B(_1479_), .Y(_1506_) );
	OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1480_), .C(index_y), .Y(_1507_) );
	AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1506_), .Y(_1508_) );
	NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1508_), .C(_1502_), .Y(_1509_) );
	NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__0_), .B(_1509__bF_buf4), .Y(_1510_) );
	OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .B(_1509__bF_buf3), .C(_1510_), .Y(_1511_) );
	NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1507_), .Y(_1512_) );
	NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_1512_), .C(_1491_), .Y(_1513_) );
	NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__0_), .B(_1513_), .Y(_1514_) );
	NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__0_), .B(_1509__bF_buf2), .Y(_1515_) );
	OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1514_), .C(_1493_), .Y(_1516_) );
	OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1511_), .C(_1516_), .Y(_1517_) );
	OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_979__bF_buf3), .C(_1123_), .Y(_1518_) );
	OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_1518_), .Y(_1519_) );
	NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1519_), .Y(_1520_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .Y(_1521_) );
	INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1522_) );
	INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .Y(_1523_) );
	NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1523_), .C(_1522_), .Y(_1524_) );
	NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1423_), .Y(_1525_) );
	NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1128_), .Y(_1526_) );
	NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1526_), .C(_1525_), .Y(_1527_) );
	NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1527_), .Y(_1528_) );
	OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1517_), .C(_1478_), .Y(AI_0_) );
	NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(ABH_1_), .B(_925__bF_buf3), .C(_1077__bF_buf2), .Y(_1529_) );
	OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1475_), .C(_1529_), .Y(_1530_) );
	AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_1_), .C(_1530_), .Y(_1531_) );
	INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .Y(_1532_) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__1_), .Y(_1533_) );
	NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .B(_1509__bF_buf1), .Y(_1534_) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__1_), .Y(_1535_) );
	NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__1_), .B(_1509__bF_buf0), .Y(_1536_) );
	OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1509__bF_buf4), .C(_1536_), .Y(_1537_) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__1_), .Y(_1538_) );
	OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1513_), .C(_1532_), .Y(_1539_) );
	OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1534_), .B(_1539_), .C(_1532_), .D(_1537_), .Y(_1540_) );
	OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1540_), .C(_1531_), .Y(AI_1_) );
	NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(ABH_2_), .B(_925__bF_buf2), .C(_1077__bF_buf1), .Y(_1541_) );
	OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_1475_), .C(_1541_), .Y(_1542_) );
	AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_2_), .C(_1542_), .Y(_1543_) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__2_), .Y(_1544_) );
	NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__2_), .B(_1509__bF_buf3), .Y(_1545_) );
	OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1509__bF_buf2), .C(_1545_), .Y(_1546_) );
	NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__2_), .B(_1513_), .Y(_1547_) );
	NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__2_), .B(_1509__bF_buf1), .Y(_1548_) );
	OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1547_), .C(_1493_), .Y(_1549_) );
	OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1546_), .C(_1549_), .Y(_1550_) );
	OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1550_), .C(_1543_), .Y(AI_2_) );
	NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(ABH_3_), .B(_925__bF_buf1), .C(_1077__bF_buf0), .Y(_1551_) );
	OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1475_), .C(_1551_), .Y(_1552_) );
	AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_3_), .C(_1552_), .Y(_1554_) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__3_), .Y(_1555_) );
	NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1509__bF_buf0), .Y(_1557_) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__3_), .Y(_1558_) );
	NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__3_), .B(_1509__bF_buf4), .Y(_1560_) );
	OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1509__bF_buf3), .C(_1560_), .Y(_1561_) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__3_), .Y(_1563_) );
	OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1513_), .C(_1532_), .Y(_1564_) );
	OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .B(_1564_), .C(_1532_), .D(_1561_), .Y(_1566_) );
	OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1566_), .C(_1554_), .Y(AI_3_) );
	INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(ABH_4_), .Y(_1568_) );
	OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_1107_), .C(_934_), .D(_1475_), .Y(_1569_) );
	AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_4_), .C(_1569_), .Y(_1571_) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__4_), .Y(_1572_) );
	NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__4_), .B(_1509__bF_buf2), .Y(_1574_) );
	OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_1509__bF_buf1), .C(_1574_), .Y(_1575_) );
	NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__4_), .B(_1513_), .Y(_1576_) );
	NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__4_), .B(_1509__bF_buf0), .Y(_1577_) );
	OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1576_), .C(_1493_), .Y(_1578_) );
	OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1575_), .C(_1578_), .Y(_84_) );
	OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_84_), .C(_1571_), .Y(AI_4_) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(ABH_5_), .Y(_85_) );
	OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_1107_), .C(_1467_), .D(_1475_), .Y(_86_) );
	AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_5_), .C(_86_), .Y(_87_) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__5_), .Y(_88_) );
	NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__5_), .B(_1509__bF_buf4), .Y(_89_) );
	OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_1509__bF_buf3), .C(_89_), .Y(_90_) );
	NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__5_), .B(_1513_), .Y(_91_) );
	NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__5_), .B(_1509__bF_buf2), .Y(_92_) );
	OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_91_), .C(_1493_), .Y(_93_) );
	OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_90_), .C(_93_), .Y(_94_) );
	OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_94_), .C(_87_), .Y(AI_5_) );
	INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(ABH_6_), .Y(_95_) );
	OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_1107_), .C(_1303_), .D(_1475_), .Y(_96_) );
	AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_6_), .C(_96_), .Y(_97_) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__6_), .Y(_98_) );
	NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__6_), .B(_1509__bF_buf1), .Y(_99_) );
	OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_1509__bF_buf0), .C(_99_), .Y(_100_) );
	NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__6_), .B(_1513_), .Y(_101_) );
	NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__6_), .B(_1509__bF_buf4), .Y(_102_) );
	OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_101_), .C(_1493_), .Y(_103_) );
	OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_100_), .C(_103_), .Y(_104_) );
	OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_104_), .C(_97_), .Y(AI_6_) );
	INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(ABH_7_), .Y(_105_) );
	OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_1107_), .C(_968_), .D(_1475_), .Y(_106_) );
	AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(ADD_7_), .C(_106_), .Y(_107_) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__7_), .Y(_108_) );
	NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_1509__bF_buf3), .Y(_109_) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__7_), .Y(_110_) );
	NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__7_), .B(_1509__bF_buf2), .Y(_112_) );
	OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_1509__bF_buf1), .C(_112_), .Y(_113_) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__7_), .Y(_115_) );
	OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_1513_), .C(_1532_), .Y(_116_) );
	OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_116_), .C(_1532_), .D(_113_), .Y(_118_) );
	OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_118_), .C(_107_), .Y(AI_7_) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(op_0_), .Y(_120_) );
	INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .Y(_121_) );
	OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_997_), .C(_925__bF_buf0), .Y(_123_) );
	NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_121_), .Y(_124_) );
	OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_121_), .C(_124_), .Y(ALU_op_0_) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(op_1_), .Y(_126_) );
	OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_121_), .C(_124_), .Y(ALU_op_1_) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(backwards), .Y(_128_) );
	OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1119_), .C(_1495_), .Y(_130_) );
	OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1094_), .C(_1236_), .Y(_131_) );
	INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
	OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf3), .B(_1104_), .C(_132_), .Y(_133_) );
	NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_133_), .Y(_134_) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
	AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(op_2_), .B(_1422_), .C(_135_), .Y(_136_) );
	OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_1107_), .C(_136_), .Y(ALU_op_2_) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(op_3_), .Y(_137_) );
	NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_121_), .Y(ALU_op_3_) );
	INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .Y(_138_) );
	NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1010_), .Y(_139_) );
	OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_979__bF_buf2), .C(_139_), .Y(_140_) );
	OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_140_), .C(store), .Y(_141_) );
	NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_141_), .C(_134_), .Y(_1603_) );
	OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1001_), .C(_134_), .Y(_142_) );
	AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(php), .Y(_143_) );
	OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_143_), .C(C), .Y(_144_) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .Y(_145_) );
	OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_1495_), .C(_1445_), .D(_132_), .Y(_146_) );
	OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(php), .B(_1523_), .C(_138_), .Y(_147_) );
	AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_147_), .C(_146_), .Y(_148_) );
	AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_144_), .Y(_149_) );
	OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_1517_), .C(_149_), .Y(_1595_) );
	INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(PC_9_), .Y(_150_) );
	NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_1540_), .Y(_151_) );
	MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(Z), .B(ADD_1_), .S(php), .Y(_152_) );
	OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_1100__bF_buf0), .C(_152_), .D(_1523_), .Y(_153_) );
	AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_1002_), .C(_153_), .Y(_154_) );
	OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_132_), .C(_154_), .Y(_155_) );
	NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_151_), .Y(_156_) );
	OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_1495_), .C(_156_), .Y(_1596_) );
	INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(PC_10_), .Y(_157_) );
	INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .Y(_158_) );
	NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(php), .B(I), .Y(_159_) );
	OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(php), .B(_158_), .C(_159_), .Y(_160_) );
	OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_1100__bF_buf3), .C(_158_), .D(_138_), .Y(_161_) );
	AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_160_), .C(_161_), .Y(_162_) );
	OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_1495_), .C(_162_), .Y(_163_) );
	AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_131_), .C(_163_), .Y(_164_) );
	OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_1550_), .C(_164_), .Y(_1597_) );
	INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(PC_11_), .Y(_165_) );
	NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_1566_), .Y(_166_) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(D), .Y(_167_) );
	MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(D), .B(ADD_3_), .S(php), .Y(_168_) );
	OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_1100__bF_buf2), .C(_168_), .D(_1523_), .Y(_169_) );
	AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_1002_), .C(_169_), .Y(_170_) );
	OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_132_), .C(_170_), .Y(_171_) );
	NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_166_), .Y(_172_) );
	OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_1495_), .C(_172_), .Y(_1598_) );
	OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_1241_), .C(ADD_4_), .D(_143_), .Y(_173_) );
	INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(PC_12_), .Y(_174_) );
	OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_1100__bF_buf1), .C(_174_), .D(_1495_), .Y(_175_) );
	AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_131_), .C(_175_), .Y(_176_) );
	AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_173_), .Y(_177_) );
	OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_84_), .C(_177_), .Y(_1599_) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(PC_13_), .Y(_178_) );
	NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_143_), .Y(_179_) );
	OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_1495_), .C(_179_), .Y(_180_) );
	OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1002_), .C(ADD_5_), .Y(_181_) );
	OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_132_), .C(_181_), .Y(_182_) );
	NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_182_), .Y(_183_) );
	OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_94_), .C(_183_), .Y(_1600_) );
	OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_143_), .C(V), .Y(_184_) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(PC_14_), .Y(_185_) );
	OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_1495_), .C(_1468_), .D(_132_), .Y(_186_) );
	AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_147_), .C(_186_), .Y(_187_) );
	AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_184_), .Y(_188_) );
	OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_104_), .C(_188_), .Y(_1601_) );
	OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_143_), .C(N), .Y(_189_) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(PC_15_), .Y(_190_) );
	OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_1495_), .C(_1469_), .D(_132_), .Y(_191_) );
	AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_147_), .C(_191_), .Y(_192_) );
	AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_189_), .Y(_193_) );
	OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_118_), .C(_193_), .Y(_1602_) );
	INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(adc_sbc), .Y(_194_) );
	NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_194_), .Y(_50_) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(adc_bcd), .Y(_195_) );
	NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_1021_), .Y(ALU_BCD) );
	INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_1257_) );
	INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(res), .Y(_198_) );
	OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_1479_), .C(_1257_), .Y(_73_) );
	NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(_1479_), .Y(_200_) );
	INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(plp), .Y(_201_) );
	OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_928__bF_buf1), .C(I), .Y(_203_) );
	OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_200_), .C(_203_), .Y(_204_) );
	NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_204_), .Y(_206_) );
	INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .Y(_207_) );
	INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(sei), .Y(_209_) );
	AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_209_), .C(cli), .Y(_210_) );
	OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_207_), .C(_1435_), .Y(_212_) );
	AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(DIMUX_2_), .C(_1095_), .Y(_213_) );
	OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_206_), .C(_213_), .Y(_27_) );
	AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(shift_right), .Y(ALU_right) );
	NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(load_reg), .B(_201_), .Y(_215_) );
	OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf0), .B(_215_), .C(_1499_), .Y(_216_) );
	OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1089_), .C(_999_), .Y(_217_) );
	NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_217_), .Y(_218_) );
	OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(RDY_bF_buf6), .Y(_219_) );
	INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(_220_) );
	NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_1513_), .Y(_221_) );
	NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_221_), .Y(_222_) );
	OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1104_), .C(ADD_0_), .Y(_223_) );
	OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1522_), .C(_223_), .Y(_224_) );
	NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_222_), .Y(_225_) );
	OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .B(_222_), .C(_225_), .Y(_1371_) );
	NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(adc_bcd), .B(adj_bcd), .C(ALU_HC), .Y(_226_) );
	NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(adj_bcd), .B(_195_), .Y(_227_) );
	OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(ALU_HC), .B(_227_), .C(_226_), .Y(_228_) );
	NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_228_), .Y(_229_) );
	INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_230_) );
	NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_230_), .Y(_231_) );
	OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_228_), .C(_231_), .Y(_232_) );
	OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1522_), .C(_232_), .Y(_233_) );
	NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_222_), .Y(_234_) );
	OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .B(_222_), .C(_234_), .Y(_1388_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(ADD_2_), .Y(_235_) );
	NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_230_), .Y(_236_) );
	NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_230_), .Y(_237_) );
	OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf4), .B(_1104_), .C(_237_), .Y(_238_) );
	OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_1522_), .C(_236_), .D(_238_), .Y(_239_) );
	NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_222_), .Y(_240_) );
	OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_222_), .C(_240_), .Y(_1395_) );
	OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_226_), .C(_237_), .Y(_241_) );
	INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .Y(_242_) );
	NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(ALU_HC), .B(_227_), .Y(_243_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_242_), .Y(_244_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_244_), .Y(_245_) );
	NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_3_), .B(_1105_), .Y(_246_) );
	OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_245_), .C(_246_), .Y(_247_) );
	NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_247_), .Y(_248_) );
	OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_222_), .C(_248_), .Y(_1402_) );
	OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1104_), .C(ADD_4_), .Y(_249_) );
	OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_1522_), .C(_249_), .Y(_250_) );
	NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_222_), .Y(_251_) );
	OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_222_), .C(_251_), .Y(_1406_) );
	INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .Y(_252_) );
	NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(adc_bcd), .C(adj_bcd), .Y(_253_) );
	INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_253_), .Y(_254_) );
	NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(_227_), .Y(_255_) );
	NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_255_), .Y(_256_) );
	NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_256_), .Y(_257_) );
	NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_256_), .Y(_258_) );
	NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_258_), .Y(_259_) );
	AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .B(_1105_), .C(_257_), .D(_259_), .Y(_260_) );
	MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_88_), .S(_222_), .Y(_1418_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(ADD_6_), .Y(_261_) );
	NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_258_), .Y(_262_) );
	OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_261_), .Y(_263_) );
	NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_262_), .C(_263_), .Y(_264_) );
	OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1522_), .C(_264_), .Y(_265_) );
	NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_222_), .Y(_266_) );
	OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_222_), .C(_266_), .Y(_1424_) );
	INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .Y(_267_) );
	OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_253_), .C(_262_), .Y(_268_) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(ADD_7_), .Y(_269_) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .Y(_270_) );
	OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1104_), .C(_270_), .Y(_271_) );
	OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_1522_), .C(_271_), .Y(_272_) );
	NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_272_), .Y(_273_) );
	OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_222_), .C(_273_), .Y(_1432_) );
	INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(NMI_1), .Y(_274_) );
	NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(NMI), .B(_937_), .C(_274_), .Y(_275_) );
	OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_1095_), .C(_275_), .Y(_28_) );
	NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(cond_code_0_), .B(_924__bF_buf2), .Y(_276_) );
	OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_1205_), .C(_276_), .Y(_58_) );
	NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_924__bF_buf0), .Y(_277_) );
	OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_1051_), .C(_277_), .Y(_59_) );
	NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(cond_code_2_), .B(_924__bF_buf6), .Y(_278_) );
	OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_1135_), .C(_278_), .Y(_60_) );
	NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf4), .B(_1143_), .Y(_279_) );
	NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_971_), .Y(_280_) );
	INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_280_), .Y(_281_) );
	NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_281_), .Y(_282_) );
	NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_282_), .Y(_283_) );
	INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_283_), .Y(_284_) );
	OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_928__bF_buf4), .C(clv), .Y(_285_) );
	OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_284_), .C(_285_), .Y(_56_) );
	NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1249_), .Y(_286_) );
	NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1143_), .Y(_287_) );
	OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_929__bF_buf3), .C(_286_), .D(_287_), .Y(_77_) );
	OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_928__bF_buf3), .C(cli), .Y(_288_) );
	OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf3), .B(_1045_), .C(_1249_), .Y(_289_) );
	OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_287_), .C(_288_), .Y(_55_) );
	OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_928__bF_buf2), .C(sed), .Y(_290_) );
	NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1051_), .Y(_291_) );
	NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_1143_), .Y(_292_) );
	OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_292_), .C(_290_), .Y(_76_) );
	OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_928__bF_buf1), .C(cld), .Y(_293_) );
	OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_292_), .C(_293_), .Y(_54_) );
	INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(sec), .Y(_294_) );
	NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1143_), .Y(_295_) );
	OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_929__bF_buf2), .C(_286_), .D(_295_), .Y(_75_) );
	OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_928__bF_buf0), .C(clc), .Y(_296_) );
	OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_295_), .C(_296_), .Y(_53_) );
	OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_928__bF_buf4), .C(php), .Y(_297_) );
	OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1301_), .B(_279_), .C(_297_), .Y(_71_) );
	OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_929__bF_buf1), .C(_1209_), .D(_279_), .Y(_72_) );
	INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(bit_ins), .Y(_298_) );
	OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf2), .B(_956_), .C(_1191_), .Y(_299_) );
	NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_1209_), .Y(_300_) );
	NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf0), .B(_300_), .Y(_301_) );
	OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_929__bF_buf4), .C(_301_), .Y(_52_) );
	NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1305_), .Y(_302_) );
	NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_302_), .C(_962_), .Y(_303_) );
	INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_303_), .Y(_304_) );
	AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_1046_), .C(_1065__bF_buf2), .Y(_305_) );
	AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_1065__bF_buf1), .C(_304_), .D(_305_), .Y(_67_) );
	OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf6), .B(_928__bF_buf3), .C(_126_), .Y(_306_) );
	NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_1038_), .Y(_307_) );
	INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_307_), .Y(_308_) );
	INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_291_), .Y(_309_) );
	NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_309_), .Y(_310_) );
	AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_1290_), .C(_1064_), .D(_308_), .Y(_311_) );
	NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_280_), .Y(_312_) );
	OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf1), .B(_1045_), .C(_951_), .Y(_313_) );
	OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_1292_), .C(_1246_), .Y(_314_) );
	AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_291_), .C(_1143_), .D(_312_), .Y(_315_) );
	INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_972_), .Y(_316_) );
	NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_1052_), .C(_1297_), .Y(_317_) );
	NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_317_), .C(_311_), .Y(_318_) );
	NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_300_), .Y(_319_) );
	OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1292_), .C(_319_), .Y(_320_) );
	NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_320_), .Y(_321_) );
	OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1292_), .C(_321_), .Y(_322_) );
	NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1292_), .Y(_323_) );
	NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf0), .B(_323_), .Y(_324_) );
	AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_1052_), .Y(_325_) );
	AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_325_), .C(_318_), .Y(_326_) );
	NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_326_), .C(_322_), .Y(_327_) );
	AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_306_), .Y(_68_) );
	OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_928__bF_buf2), .C(op_2_), .Y(_328_) );
	OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf3), .B(_321_), .C(_328_), .Y(_69_) );
	AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_1065__bF_buf2), .C(_324_), .D(_319_), .Y(_70_) );
	INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_329_) );
	NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .Y(_330_) );
	INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(_330_), .Y(_331_) );
	OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__0_), .Y(_332_) );
	OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_331_), .C(_332_), .Y(_1553_) );
	INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(_333_) );
	OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__1_), .Y(_334_) );
	OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_331_), .C(_334_), .Y(_1556_) );
	INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_335_) );
	OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__2_), .Y(_336_) );
	OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_331_), .C(_336_), .Y(_1559_) );
	INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_247_), .Y(_337_) );
	OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__3_), .Y(_338_) );
	OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_337_), .C(_338_), .Y(_1562_) );
	INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_250_), .Y(_339_) );
	OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__4_), .Y(_340_) );
	OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_331_), .C(_340_), .Y(_1565_) );
	OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__5_), .Y(_341_) );
	OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_331_), .C(_341_), .Y(_1567_) );
	INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_265_), .Y(_342_) );
	OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__6_), .Y(_343_) );
	OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_331_), .C(_343_), .Y(_1570_) );
	INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_272_), .Y(_344_) );
	OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_221_), .C(AXYS_2__7_), .Y(_345_) );
	OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_344_), .C(_345_), .Y(_1573_) );
	NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1205_), .Y(_346_) );
	NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_1046_), .Y(_347_) );
	NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_1292_), .Y(_348_) );
	AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_1135_), .C(_346_), .D(_1297_), .Y(_349_) );
	OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_928__bF_buf1), .C(rotate), .Y(_350_) );
	OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf1), .B(_349_), .C(_350_), .Y(_74_) );
	NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1306_), .Y(_351_) );
	INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_351_), .Y(_352_) );
	OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_928__bF_buf0), .C(shift_right), .Y(_353_) );
	OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf0), .B(_352_), .C(_353_), .Y(_79_) );
	AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_971_), .C(_1065__bF_buf3), .Y(_354_) );
	AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1065__bF_buf2), .C(_311_), .D(_354_), .Y(_57_) );
	NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf3), .B(_1278_), .C(_323_), .Y(_355_) );
	OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_929__bF_buf2), .C(_355_), .Y(_78_) );
	OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1167_), .C(_925__bF_buf5), .Y(_356_) );
	NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_356_), .Y(_357_) );
	NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(D), .B(_1135_), .Y(_358_) );
	NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_302_), .Y(_359_) );
	NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_359_), .Y(_360_) );
	OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_357_), .C(_358_), .D(_360_), .Y(_48_) );
	OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_357_), .C(_360_), .Y(_49_) );
	AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_348_), .C(_1143_), .D(_310_), .Y(_361_) );
	OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_928__bF_buf4), .C(inc), .Y(_362_) );
	OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf1), .B(_361_), .C(_362_), .Y(_63_) );
	OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_928__bF_buf3), .C(load_only), .Y(_363_) );
	OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf0), .B(_282_), .C(_363_), .Y(_65_) );
	INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .Y(_364_) );
	NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_1067_), .C(_364_), .Y(_365_) );
	OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_929__bF_buf1), .C(_365_), .Y(_83_) );
	NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_1509__bF_buf0), .Y(_366_) );
	NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_366_), .Y(_367_) );
	NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__0_), .B(_367_), .Y(_368_) );
	AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_367_), .C(_368_), .Y(_111_) );
	NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_367_), .Y(_369_) );
	OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_367_), .C(_369_), .Y(_114_) );
	NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__2_), .B(_367_), .Y(_370_) );
	AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_367_), .C(_370_), .Y(_117_) );
	NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_247_), .Y(_371_) );
	OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_367_), .C(_371_), .Y(_119_) );
	NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__4_), .B(_367_), .Y(_372_) );
	AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_367_), .C(_372_), .Y(_122_) );
	NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__5_), .B(_367_), .Y(_373_) );
	AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_367_), .C(_373_), .Y(_125_) );
	NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__6_), .B(_367_), .Y(_374_) );
	AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_367_), .C(_374_), .Y(_127_) );
	NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_272_), .Y(_375_) );
	OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_367_), .C(_375_), .Y(_129_) );
	NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_280_), .Y(_376_) );
	OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_1191_), .C(_376_), .Y(_377_) );
	OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf7), .B(_928__bF_buf2), .C(store), .Y(_378_) );
	OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1065__bF_buf3), .B(_377_), .C(_378_), .Y(_82_) );
	OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf6), .B(_928__bF_buf1), .C(index_y), .Y(_379_) );
	OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1232_), .C(_929__bF_buf0), .Y(_380_) );
	NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_1292_), .Y(_381_) );
	NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1067_), .C(_381_), .Y(_382_) );
	NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_382_), .C(_380_), .Y(_64_) );
	INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(src_reg_0_), .Y(_383_) );
	INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .Y(_384_) );
	NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1143_), .Y(_385_) );
	OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf0), .B(_1045_), .C(_971_), .Y(_386_) );
	OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_386_), .Y(_387_) );
	OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_307_), .C(_387_), .Y(_388_) );
	NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_376_), .Y(_389_) );
	INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_313_), .Y(_390_) );
	NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_281_), .C(_390_), .Y(_391_) );
	OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_389_), .C(_391_), .Y(_392_) );
	NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_388_), .Y(_393_) );
	OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_284_), .C(_393_), .Y(_394_) );
	NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_929__bF_buf4), .B(_394_), .Y(_395_) );
	OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_929__bF_buf3), .C(_395_), .Y(_80_) );
	INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(src_reg_1_), .Y(_396_) );
	NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1297_), .Y(_397_) );
	OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_397_), .C(_929__bF_buf2), .Y(_398_) );
	NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_947_), .Y(_399_) );
	OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_399_), .C(_381_), .Y(_400_) );
	OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_307_), .C(_400_), .Y(_401_) );
	NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_398_), .Y(_402_) );
	AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_1065__bF_buf2), .C(_402_), .D(_393_), .Y(_81_) );
	INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_0_), .Y(_403_) );
	OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_951_), .C(_1038_), .Y(_404_) );
	OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_404_), .C(_387_), .Y(_405_) );
	OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_384_), .C(_1273_), .Y(_406_) );
	OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_405_), .C(_929__bF_buf1), .Y(_407_) );
	OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_929__bF_buf0), .C(_407_), .Y(_61_) );
	INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_1_), .Y(_408_) );
	INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_405_), .Y(_409_) );
	OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_282_), .C(_1184_), .D(_292_), .Y(_410_) );
	NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_410_), .Y(_411_) );
	AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_1065__bF_buf1), .C(_411_), .D(_409_), .Y(_62_) );
	INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(load_reg), .Y(_412_) );
	NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_283_), .Y(_413_) );
	NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1051_), .C(_973_), .Y(_414_) );
	OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf4), .B(_960_), .C(_1066_), .Y(_415_) );
	NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_280_), .Y(_416_) );
	AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_416_), .C(_1042_), .D(_1297_), .Y(_417_) );
	NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_417_), .C(_413_), .Y(_418_) );
	NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .B(_283_), .Y(_419_) );
	NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_309_), .Y(_420_) );
	AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_386_), .C(_1297_), .D(_420_), .Y(_421_) );
	NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_421_), .C(_419_), .Y(_422_) );
	OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .C(_929__bF_buf4), .Y(_423_) );
	OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_929__bF_buf3), .C(_423_), .Y(_66_) );
	NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1257_), .C(_1518_), .Y(_424_) );
	OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf5), .B(_928__bF_buf0), .C(IRHOLD_valid), .Y(_425_) );
	OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_425_), .C(_424_), .Y(_26_) );
	NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_366_), .Y(_426_) );
	NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__0_), .B(_426_), .Y(_427_) );
	AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_426_), .C(_427_), .Y(_196_) );
	NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__1_), .B(_426_), .Y(_428_) );
	AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_426_), .C(_428_), .Y(_197_) );
	NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__2_), .B(_426_), .Y(_429_) );
	AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_426_), .C(_429_), .Y(_199_) );
	NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__3_), .B(_426_), .Y(_430_) );
	AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_426_), .C(_430_), .Y(_202_) );
	NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__4_), .B(_426_), .Y(_431_) );
	AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_426_), .C(_431_), .Y(_205_) );
	NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__5_), .B(_426_), .Y(_432_) );
	AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_426_), .C(_432_), .Y(_208_) );
	NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__6_), .B(_426_), .Y(_433_) );
	AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_426_), .C(_433_), .Y(_211_) );
	NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__7_), .B(_426_), .Y(_434_) );
	AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_426_), .C(_434_), .Y(_214_) );
	NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_0_), .B(_424_), .Y(_435_) );
	OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_424_), .C(_435_), .Y(_18_) );
	NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_1_), .B(_424_), .Y(_436_) );
	OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_424_), .C(_436_), .Y(_19_) );
	NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_2_), .B(_424_), .Y(_437_) );
	OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_424_), .C(_437_), .Y(_20_) );
	NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_3_), .B(_424_), .Y(_438_) );
	OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_424_), .C(_438_), .Y(_21_) );
	MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_934_), .S(_424_), .Y(_22_) );
	INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_5_), .Y(_439_) );
	MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_1467_), .S(_424_), .Y(_23_) );
	MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1303_), .S(_424_), .Y(_24_) );
	INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_7_), .Y(_440_) );
	MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_968_), .S(_424_), .Y(_25_) );
	NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_1021_), .Y(_441_) );
	OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_441_), .C(DIMUX_6_), .Y(_442_) );
	INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_441_), .Y(_443_) );
	AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_194_), .C(plp), .Y(_444_) );
	OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(ALU_V), .C(_444_), .Y(_445_) );
	OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_201_), .C(clv), .D(_445_), .Y(_446_) );
	NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_1479_), .Y(_447_) );
	AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_446_), .C(_447_), .D(_443_), .Y(_448_) );
	OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_448_), .C(_442_), .Y(_46_) );
	NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(cld), .Y(_449_) );
	OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(D), .B(sed), .C(_449_), .Y(_450_) );
	OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_201_), .C(_450_), .Y(_451_) );
	OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_1479_), .C(_1435_), .Y(_452_) );
	AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_451_), .C(_452_), .Y(_453_) );
	AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1081_), .C(_453_), .Y(_17_) );
	NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(ALU_N), .B(_1002_), .Y(_454_) );
	INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .Y(_455_) );
	NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_1502_), .Y(_456_) );
	NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_456_), .C(_1509__bF_buf4), .Y(_457_) );
	AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(load_reg), .C(compare), .Y(_458_) );
	NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(N), .B(_458_), .Y(_459_) );
	OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1513_), .C(load_reg), .Y(_460_) );
	NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_460_), .Y(_461_) );
	AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(ALU_N), .C(plp), .Y(_462_) );
	NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_462_), .Y(_463_) );
	INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .Y(_464_) );
	AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(plp), .C(_928__bF_buf4), .Y(_465_) );
	NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_441_), .Y(_466_) );
	OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(N), .B(_441_), .C(_466_), .Y(_467_) );
	OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_467_), .C(_1435_), .Y(_468_) );
	AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_465_), .C(_468_), .Y(_469_) );
	OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_7_), .B(_1435_), .C(_138_), .Y(_470_) );
	OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_469_), .C(_454_), .Y(_29_) );
	NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(ALU_Z), .B(_1002_), .Y(_471_) );
	NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_298_), .C(_460_), .Y(_472_) );
	NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(ALU_Z), .B(_472_), .Y(_473_) );
	NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(Z), .B(_298_), .C(_458_), .Y(_474_) );
	NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_473_), .C(_474_), .Y(_475_) );
	INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .Y(_476_) );
	AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(plp), .C(_928__bF_buf3), .Y(_477_) );
	OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_1479_), .C(_1435_), .Y(_478_) );
	AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_478_), .Y(_479_) );
	OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .B(_1435_), .C(_138_), .Y(_480_) );
	OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_479_), .C(_471_), .Y(_47_) );
	INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .Y(_481_) );
	NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(shift), .B(_1002_), .Y(_482_) );
	NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(write_back), .B(_928__bF_buf2), .Y(_483_) );
	NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1427_), .C(_194_), .Y(_484_) );
	NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_294_), .Y(_485_) );
	NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(clc), .Y(_486_) );
	AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(plp), .C(_486_), .D(_485_), .Y(_487_) );
	NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(_484_), .Y(_488_) );
	OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_487_), .C(_488_), .Y(_489_) );
	OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_483_), .C(_1435_), .Y(_490_) );
	AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_483_), .C(_490_), .Y(_491_) );
	OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(_1435_), .C(_482_), .Y(_492_) );
	OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_482_), .C(_492_), .D(_491_), .Y(_16_) );
	NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(DI_7_), .Y(_493_) );
	OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_128_), .C(_493_), .Y(_51_) );
	OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1005__bF_buf1), .C(_1435_), .Y(_494_) );
	AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_1086_), .C(_494_), .Y(_495_) );
	NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .B(_1500_), .C(_495_), .Y(_496_) );
	OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_999_), .C(_1235_), .Y(_497_) );
	OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_979__bF_buf1), .C(_497_), .Y(_498_) );
	AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf4), .B(_1027_), .C(_1075_), .Y(_499_) );
	OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1005__bF_buf0), .C(_499_), .Y(_500_) );
	NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_500_), .Y(_501_) );
	NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1071_), .Y(_502_) );
	OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf0), .B(_988_), .C(_502_), .Y(_503_) );
	NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_503_), .Y(_504_) );
	NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_501_), .Y(_505_) );
	NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_505_), .Y(_506_) );
	OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001_), .C(_1421_), .Y(_507_) );
	OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_1267_), .Y(_508_) );
	NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(_130_), .Y(_509_) );
	NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .B(_1010_), .Y(_510_) );
	OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf2), .B(_1252_), .C(_510_), .Y(_511_) );
	OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf4), .B(_1119_), .C(_994_), .Y(_512_) );
	NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_511_), .Y(_513_) );
	NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_513_), .Y(_514_) );
	NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_514_), .Y(_515_) );
	NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_515_), .Y(_516_) );
	INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_517_) );
	AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(ABH_0_), .C(ADD_0_), .D(_511_), .Y(_518_) );
	NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_509_), .C(_518_), .Y(_519_) );
	OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_496_), .Y(_520_) );
	AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(_517_), .C(_520_), .Y(_521_) );
	OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_516_), .C(_521_), .Y(_1593_) );
	INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(ABH_0_), .Y(_522_) );
	OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1086_), .C(_1006_), .Y(_523_) );
	NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_499_), .C(_510_), .Y(_524_) );
	NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_1020_), .Y(_525_) );
	NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_1007_), .C(_992_), .Y(_526_) );
	OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_526_), .C(_990_), .Y(_527_) );
	NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_525_), .Y(_528_) );
	INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_528_), .Y(_529_) );
	NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .B(_502_), .C(_529_), .Y(_530_) );
	NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_530_), .Y(_531_) );
	NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1237_), .Y(_532_) );
	AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_1258_), .C(_1171_), .Y(_533_) );
	NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_532_), .C(_1263_), .Y(_534_) );
	NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1163_), .Y(_535_) );
	NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1325_), .Y(_536_) );
	NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .Y(_537_) );
	AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_1015_), .C(_1431_), .Y(_538_) );
	OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_1162_), .C(_538_), .Y(_539_) );
	OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_537_), .Y(_540_) );
	NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_540_), .Y(_541_) );
	AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_1496_), .C(_999_), .D(_1077__bF_buf3), .Y(_542_) );
	OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf3), .B(_980__bF_buf1), .C(_542_), .Y(_543_) );
	OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_1009_), .C(_497_), .Y(_544_) );
	OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf2), .B(_925__bF_buf3), .C(_1236_), .Y(_545_) );
	NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_544_), .Y(_546_) );
	AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1077__bF_buf2), .B(_998_), .C(_1006_), .D(_1089_), .Y(_547_) );
	NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_546_), .Y(_548_) );
	NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_548_), .Y(_549_) );
	NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_542_), .C(_547_), .Y(_550_) );
	OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf1), .B(_990_), .C(_1236_), .Y(_551_) );
	OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_551_), .Y(_552_) );
	NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_552_), .Y(_553_) );
	OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_549_), .C(_541_), .Y(_554_) );
	OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1154_), .C(_533_), .Y(_555_) );
	INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .Y(_556_) );
	NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1431_), .Y(_557_) );
	NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_356_), .C(_557_), .Y(_558_) );
	INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .Y(_559_) );
	NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1241_), .Y(_560_) );
	NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_1526_), .C(_560_), .Y(_561_) );
	OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_555_), .C(_561_), .D(_558_), .Y(_562_) );
	NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1450_), .Y(_563_) );
	NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1448_), .C(_563_), .Y(_564_) );
	OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_543_), .Y(_565_) );
	NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_565_), .Y(_566_) );
	NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_562_), .C(_566_), .Y(_567_) );
	NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_554_), .Y(_568_) );
	OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_528_), .Y(_569_) );
	OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_550_), .Y(_570_) );
	OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_979__bF_buf0), .B(_1000__bF_buf2), .C(_1236_), .Y(_571_) );
	OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_979__bF_buf3), .C(_1096_), .Y(_572_) );
	OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_571_), .Y(_573_) );
	OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_503_), .Y(_574_) );
	NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_574_), .Y(_575_) );
	NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_575_), .Y(_576_) );
	OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_576_), .C(RDY_bF_buf2), .Y(_577_) );
	AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_531_), .C(_577_), .Y(_578_) );
	NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_578__bF_buf4), .Y(_579_) );
	OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_578__bF_buf3), .C(_579_), .Y(_0_) );
	INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(_511_), .Y(_580_) );
	OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_507_), .C(ABH_1_), .Y(_581_) );
	OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_580_), .C(_581_), .Y(_582_) );
	AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .B(_517_), .C(_582_), .Y(_583_) );
	OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_516_), .C(_583_), .Y(_1594_) );
	INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(ABH_1_), .Y(_584_) );
	NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(_578__bF_buf2), .Y(_585_) );
	OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_578__bF_buf1), .C(_585_), .Y(_1_) );
	OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_580_), .C(_948_), .D(_501_), .Y(_586_) );
	AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(ABH_2_), .B(_508_), .C(_586_), .Y(_587_) );
	OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_516_), .C(_587_), .Y(_1580_) );
	INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(ABH_2_), .Y(_588_) );
	NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_578__bF_buf0), .Y(_589_) );
	OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_578__bF_buf4), .C(_589_), .Y(_2_) );
	OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_580_), .C(_1138_), .D(_501_), .Y(_590_) );
	AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(ABH_3_), .B(_508_), .C(_590_), .Y(_591_) );
	OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_516_), .C(_591_), .Y(_1581_) );
	INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(ABH_3_), .Y(_592_) );
	NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_578__bF_buf3), .Y(_593_) );
	OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_578__bF_buf2), .C(_593_), .Y(_3_) );
	INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .Y(_594_) );
	OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_580_), .C(_934_), .D(_501_), .Y(_595_) );
	AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(ABH_4_), .B(_508_), .C(_595_), .Y(_596_) );
	OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_516_), .C(_596_), .Y(_1582_) );
	NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_578__bF_buf1), .Y(_597_) );
	OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_578__bF_buf0), .C(_597_), .Y(_4_) );
	OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_507_), .C(ABH_5_), .Y(_598_) );
	OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_580_), .C(_598_), .Y(_599_) );
	AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .B(_517_), .C(_599_), .Y(_600_) );
	OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_516_), .C(_600_), .Y(_1583_) );
	NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .B(_578__bF_buf4), .Y(_601_) );
	OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_578__bF_buf3), .C(_601_), .Y(_5_) );
	OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_580_), .C(_1303_), .D(_501_), .Y(_602_) );
	AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(ABH_6_), .B(_508_), .C(_602_), .Y(_603_) );
	OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_516_), .C(_603_), .Y(_1584_) );
	NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1584_), .B(_578__bF_buf2), .Y(_604_) );
	OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_578__bF_buf1), .C(_604_), .Y(_6_) );
	OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_507_), .C(ABH_7_), .Y(_605_) );
	OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_580_), .C(_605_), .Y(_606_) );
	AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_7_), .B(_517_), .C(_606_), .Y(_607_) );
	OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_516_), .C(_607_), .Y(_1585_) );
	NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_578__bF_buf0), .Y(_608_) );
	OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_578__bF_buf4), .C(_608_), .Y(_7_) );
	NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_1517_), .Y(_609_) );
	INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(_506_), .Y(_610_) );
	INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(ABL_0_), .Y(_611_) );
	AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_1267_), .C(DIMUX_0_), .D(_512_), .Y(_612_) );
	NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_511_), .Y(_613_) );
	OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
	AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_0_), .C(_614_), .Y(_615_) );
	OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_516_), .C(_615_), .Y(_616_) );
	OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_609_), .Y(_1579_) );
	OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_616_), .C(_578__bF_buf3), .Y(_617_) );
	OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_578__bF_buf2), .C(_617_), .Y(_8_) );
	NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_1540_), .Y(_618_) );
	INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(ABL_1_), .Y(_619_) );
	AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_1_), .C(DIMUX_1_), .D(_512_), .Y(_620_) );
	OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_613_), .C(_620_), .Y(_621_) );
	AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_1_), .C(_621_), .Y(_622_) );
	OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_516_), .C(_622_), .Y(_623_) );
	OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_618_), .Y(_1586_) );
	OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_623_), .C(_578__bF_buf1), .Y(_624_) );
	OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_578__bF_buf0), .C(_624_), .Y(_9_) );
	NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_1550_), .Y(_625_) );
	INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(ABL_2_), .Y(_626_) );
	AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_2_), .C(DIMUX_2_), .D(_512_), .Y(_627_) );
	OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_613_), .C(_627_), .Y(_628_) );
	AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_2_), .C(_628_), .Y(_629_) );
	OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_516_), .C(_629_), .Y(_630_) );
	OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_625_), .Y(_1587_) );
	OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_630_), .C(_578__bF_buf4), .Y(_631_) );
	OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_578__bF_buf3), .C(_631_), .Y(_10_) );
	NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_1566_), .Y(_632_) );
	INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(ABL_3_), .Y(_633_) );
	AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_3_), .C(DIMUX_3_), .D(_512_), .Y(_634_) );
	OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_613_), .C(_634_), .Y(_635_) );
	AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_3_), .C(_635_), .Y(_636_) );
	OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_516_), .C(_636_), .Y(_637_) );
	OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(_632_), .Y(_1588_) );
	OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_637_), .C(_578__bF_buf2), .Y(_638_) );
	OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_578__bF_buf1), .C(_638_), .Y(_11_) );
	NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_84_), .Y(_639_) );
	INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(ABL_4_), .Y(_640_) );
	AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_4_), .C(DIMUX_4_), .D(_512_), .Y(_641_) );
	OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_613_), .C(_641_), .Y(_642_) );
	AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_4_), .C(_642_), .Y(_643_) );
	OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_516_), .C(_643_), .Y(_644_) );
	OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_639_), .Y(_1589_) );
	OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_644_), .C(_578__bF_buf0), .Y(_645_) );
	OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_578__bF_buf4), .C(_645_), .Y(_12_) );
	NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_94_), .Y(_646_) );
	INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(ABL_5_), .Y(_647_) );
	AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_5_), .C(DIMUX_5_), .D(_512_), .Y(_648_) );
	OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_613_), .C(_648_), .Y(_649_) );
	AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_5_), .C(_649_), .Y(_650_) );
	OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_516_), .C(_650_), .Y(_651_) );
	OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_646_), .Y(_1590_) );
	OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_651_), .C(_578__bF_buf3), .Y(_652_) );
	OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_578__bF_buf2), .C(_652_), .Y(_13_) );
	NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_104_), .Y(_653_) );
	INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(ABL_6_), .Y(_654_) );
	AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_6_), .C(DIMUX_6_), .D(_512_), .Y(_655_) );
	OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_613_), .C(_655_), .Y(_656_) );
	AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_6_), .C(_656_), .Y(_657_) );
	OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_516_), .C(_657_), .Y(_658_) );
	OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_653_), .Y(_1591_) );
	OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_658_), .C(_578__bF_buf1), .Y(_659_) );
	OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_578__bF_buf0), .C(_659_), .Y(_14_) );
	NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_118_), .Y(_660_) );
	INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(ABL_7_), .Y(_661_) );
	AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ADD_7_), .C(DIMUX_7_), .D(_512_), .Y(_662_) );
	OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_613_), .C(_662_), .Y(_663_) );
	AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(ADD_7_), .C(_663_), .Y(_664_) );
	OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_516_), .C(_664_), .Y(_665_) );
	OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_660_), .Y(_1592_) );
	OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_665_), .C(_578__bF_buf4), .Y(_666_) );
	OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_578__bF_buf3), .C(_666_), .Y(_15_) );
	AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1005__bF_buf3), .Y(_667_) );
	NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_667_), .Y(_668_) );
	OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1074_), .C(_1014_), .D(_667_), .Y(_669_) );
	NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .Y(_670_) );
	OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1089_), .C(_925__bF_buf2), .Y(_671_) );
	OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_1077__bF_buf1), .C(_925__bF_buf1), .Y(_672_) );
	AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_672_), .Y(_673_) );
	NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_673_), .Y(_674_) );
	AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_999_), .C(_1004_), .D(_1006_), .Y(_675_) );
	OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_1160_), .C(_675_), .Y(_676_) );
	NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_925__bF_buf0), .C(_1077__bF_buf0), .Y(_677_) );
	NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(PC_0_), .B(_925__bF_buf5), .C(_526_), .Y(_678_) );
	NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(ABL_0_), .B(_953__bF_buf3), .Y(_679_) );
	OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_953__bF_buf2), .C(_679_), .Y(_680_) );
	NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_680_), .Y(_681_) );
	NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_678_), .C(_681_), .Y(_682_) );
	AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_676_), .C(_682_), .Y(_683_) );
	OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_674_), .C(_683_), .Y(_684_) );
	NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_953__bF_buf1), .B(_928__bF_buf1), .Y(_685_) );
	OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_1108_), .C(_497_), .Y(_686_) );
	NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_686_), .Y(_687_) );
	OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf0), .B(_1094_), .C(_1170_), .Y(_688_) );
	OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_1074_), .C(state_4_), .D(_1014_), .Y(_689_) );
	NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_689_), .Y(_690_) );
	OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_980__bF_buf4), .B(_1119_), .C(_1146_), .Y(_691_) );
	INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_691_), .Y(_692_) );
	NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_692_), .C(_687_), .Y(_693_) );
	NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_684_), .Y(_694_) );
	NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_672_), .Y(_695_) );
	NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_676_), .C(_695_), .Y(_696_) );
	OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(ADD_0_), .Y(_697_) );
	AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_678_), .Y(_698_) );
	NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_698_), .C(_697_), .Y(_699_) );
	OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_696_), .C(_693_), .Y(_700_) );
	NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_700_), .Y(_701_) );
	OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1445_), .C(_701_), .D(_694_), .Y(_30_) );
	NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(PC_0_), .B(_670_), .C(_673_), .Y(_702_) );
	AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_692_), .Y(_703_) );
	AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_703_), .C(_702_), .D(_683_), .Y(_704_) );
	NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_1111_), .Y(_705_) );
	OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_695_), .C(_705_), .Y(_706_) );
	INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_706_), .Y(_707_) );
	NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf0), .B(_939__bF_buf0), .Y(_708_) );
	OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_1107_), .C(res), .D(_1100__bF_buf0), .Y(_709_) );
	AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(ABL_1_), .B(_708_), .C(_709_), .Y(_710_) );
	OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_670_), .C(_710_), .Y(_711_) );
	INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_711_), .Y(_712_) );
	OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_707_), .C(_712_), .Y(_713_) );
	NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_713_), .Y(_714_) );
	AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(PC_1_), .C(_711_), .Y(_715_) );
	OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_700_), .C(RDY_bF_buf8), .Y(_716_) );
	OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1461_), .C(_716_), .D(_714_), .Y(_37_) );
	NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_700_), .Y(_717_) );
	AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_158_), .Y(_718_) );
	NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_925__bF_buf4), .C(_1077__bF_buf3), .Y(_719_) );
	NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(res), .B(_937_), .Y(_720_) );
	INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_720_), .Y(_721_) );
	NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf3), .B(_721_), .C(_1089_), .Y(_722_) );
	NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_925__bF_buf2), .C(_526_), .Y(_723_) );
	NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_719_), .C(_722_), .Y(_724_) );
	NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(ABL_2_), .B(_953__bF_buf0), .Y(_725_) );
	OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_953__bF_buf4), .C(_725_), .Y(_726_) );
	AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_1479_), .Y(_727_) );
	NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_718_), .C(_727_), .Y(_728_) );
	OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_674_), .C(_728_), .Y(_729_) );
	NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_717_), .Y(_730_) );
	NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_676_), .C(_695_), .Y(_731_) );
	OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(ADD_2_), .Y(_732_) );
	OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_1107_), .C(_1100__bF_buf3), .D(_720_), .Y(_733_) );
	AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_1111_), .C(_733_), .Y(_734_) );
	NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_726_), .Y(_735_) );
	NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_734_), .C(_732_), .Y(_736_) );
	OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_736_), .C(_717_), .Y(_737_) );
	NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_737_), .Y(_738_) );
	OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1463_), .C(_730_), .D(_738_), .Y(_38_) );
	AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_242_), .Y(_739_) );
	NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_925__bF_buf1), .C(_1077__bF_buf2), .Y(_740_) );
	NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_925__bF_buf0), .C(_526_), .Y(_741_) );
	NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf2), .B(_741_), .C(_740_), .Y(_742_) );
	NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_939__bF_buf3), .Y(_743_) );
	NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(ABL_3_), .B(_953__bF_buf3), .Y(_744_) );
	AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_744_), .C(_928__bF_buf4), .Y(_745_) );
	NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_742_), .C(_739_), .Y(_746_) );
	OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_674_), .C(_746_), .Y(_747_) );
	AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_729_), .C(_747_), .Y(_748_) );
	NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_670_), .C(_673_), .Y(_749_) );
	NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_670_), .C(_673_), .Y(_750_) );
	AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_750_), .C(_749_), .D(_728_), .Y(_751_) );
	NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_704_), .C(_713_), .Y(_752_) );
	NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_752_), .Y(_753_) );
	OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1464_), .C(_753_), .D(_748_), .Y(_39_) );
	NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_676_), .C(_695_), .Y(_754_) );
	OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(ADD_3_), .Y(_755_) );
	OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_1107_), .C(_1100__bF_buf1), .Y(_756_) );
	AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_1111_), .C(_756_), .Y(_757_) );
	OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_953__bF_buf2), .C(_744_), .Y(_758_) );
	NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_758_), .Y(_759_) );
	NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_757_), .C(_755_), .Y(_760_) );
	OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_760_), .C(_731_), .D(_736_), .Y(_761_) );
	NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_700_), .C(_761_), .Y(_762_) );
	AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_594_), .Y(_763_) );
	NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_925__bF_buf5), .C(_1077__bF_buf1), .Y(_764_) );
	NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_925__bF_buf4), .C(_526_), .Y(_765_) );
	NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf0), .B(_765_), .C(_764_), .Y(_766_) );
	NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_939__bF_buf2), .Y(_767_) );
	NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(ABL_4_), .B(_953__bF_buf1), .Y(_768_) );
	AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_768_), .C(_928__bF_buf3), .Y(_769_) );
	NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_766_), .C(_763_), .Y(_770_) );
	OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_674_), .C(_770_), .Y(_771_) );
	NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_762_), .Y(_772_) );
	INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_771_), .Y(_773_) );
	OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_752_), .C(RDY_bF_buf2), .Y(_774_) );
	OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1465_), .C(_774_), .D(_772_), .Y(_40_) );
	AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_252_), .Y(_775_) );
	NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .B(_925__bF_buf3), .C(_1077__bF_buf0), .Y(_776_) );
	NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_925__bF_buf2), .C(_526_), .Y(_777_) );
	NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf3), .B(_777_), .C(_776_), .Y(_778_) );
	NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_939__bF_buf1), .Y(_779_) );
	NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(ABL_5_), .B(_953__bF_buf0), .Y(_780_) );
	AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_780_), .C(_928__bF_buf2), .Y(_781_) );
	NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_778_), .C(_775_), .Y(_782_) );
	OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_674_), .C(_782_), .Y(_783_) );
	AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_771_), .C(_783_), .Y(_784_) );
	NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_670_), .C(_673_), .Y(_785_) );
	NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_670_), .C(_673_), .Y(_786_) );
	AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_785_), .C(_786_), .D(_782_), .Y(_787_) );
	INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_787_), .Y(_788_) );
	OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_752_), .C(RDY_bF_buf0), .Y(_789_) );
	OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1466_), .C(_789_), .D(_784_), .Y(_41_) );
	AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_267_), .Y(_790_) );
	NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_925__bF_buf1), .C(_1077__bF_buf3), .Y(_791_) );
	NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .B(_925__bF_buf0), .C(_526_), .Y(_792_) );
	NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf2), .B(_792_), .C(_791_), .Y(_793_) );
	NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .B(_939__bF_buf0), .Y(_794_) );
	NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(ABL_6_), .B(_953__bF_buf4), .Y(_795_) );
	AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_795_), .C(_928__bF_buf1), .Y(_796_) );
	NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_793_), .C(_790_), .Y(_797_) );
	OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_674_), .C(_797_), .Y(_798_) );
	AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_787_), .C(_798_), .Y(_799_) );
	NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_798_), .C(_762_), .Y(_800_) );
	NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_800_), .Y(_801_) );
	OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1468_), .C(_799_), .D(_801_), .Y(_42_) );
	AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_464_), .Y(_802_) );
	NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_925__bF_buf5), .C(_1077__bF_buf2), .Y(_803_) );
	NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .B(_925__bF_buf4), .C(_526_), .Y(_804_) );
	NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf1), .B(_804_), .C(_803_), .Y(_805_) );
	MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(ABL_7_), .B(PC_7_), .S(_953__bF_buf3), .Y(_806_) );
	NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf0), .B(_806_), .Y(_807_) );
	NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_807_), .C(_802_), .Y(_808_) );
	OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_674_), .C(_808_), .Y(_809_) );
	INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_810_) );
	AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_810_), .Y(_811_) );
	NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .B(_670_), .C(_673_), .Y(_812_) );
	NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .B(_670_), .C(_673_), .Y(_813_) );
	AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_812_), .C(_813_), .D(_808_), .Y(_814_) );
	NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_814_), .Y(_815_) );
	OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_752_), .C(RDY_bF_buf5), .Y(_816_) );
	OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1469_), .C(_816_), .D(_811_), .Y(_43_) );
	NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .B(_924__bF_buf4), .Y(_817_) );
	NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_752_), .Y(_818_) );
	AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_1446_), .Y(_819_) );
	NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_925__bF_buf3), .C(_526_), .Y(_820_) );
	NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf0), .B(_820_), .C(_1476_), .Y(_821_) );
	NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .B(_939__bF_buf3), .Y(_822_) );
	NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(ABH_0_), .B(_953__bF_buf2), .Y(_823_) );
	AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_823_), .C(_928__bF_buf4), .Y(_824_) );
	NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_821_), .C(_819_), .Y(_825_) );
	OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_674_), .C(_825_), .Y(_826_) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_826_), .Y(_827_) );
	OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_827_), .C(_817_), .Y(_44_) );
	AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_1462_), .Y(_828_) );
	NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_925__bF_buf2), .C(_526_), .Y(_829_) );
	NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf3), .B(_829_), .C(_1529_), .Y(_830_) );
	MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(ABH_1_), .B(PC_9_), .S(_953__bF_buf1), .Y(_831_) );
	NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf3), .B(_831_), .Y(_832_) );
	NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_832_), .C(_828_), .Y(_833_) );
	OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_674_), .C(_833_), .Y(_834_) );
	AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_826_), .C(_834_), .Y(_835_) );
	AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_814_), .Y(_836_) );
	NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .B(_670_), .C(_673_), .Y(_837_) );
	NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(PC_9_), .B(_670_), .C(_673_), .Y(_838_) );
	AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_837_), .C(_838_), .D(_833_), .Y(_839_) );
	NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_839_), .C(_762_), .Y(_840_) );
	NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_840_), .Y(_841_) );
	OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_150_), .C(_841_), .D(_835_), .Y(_45_) );
	INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_840_), .Y(_842_) );
	AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_948_), .Y(_843_) );
	NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_925__bF_buf1), .C(_526_), .Y(_844_) );
	NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf2), .B(_844_), .C(_1541_), .Y(_845_) );
	NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(PC_10_), .B(_939__bF_buf2), .Y(_846_) );
	NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(ABH_2_), .B(_953__bF_buf0), .Y(_847_) );
	AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_847_), .C(_928__bF_buf2), .Y(_848_) );
	NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_845_), .C(_843_), .Y(_849_) );
	OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_674_), .C(_849_), .Y(_850_) );
	NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_842_), .Y(_851_) );
	INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_850_), .Y(_852_) );
	OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_840_), .C(RDY_bF_buf1), .Y(_853_) );
	OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_157_), .C(_853_), .D(_851_), .Y(_31_) );
	AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_497_), .C(_1138_), .Y(_854_) );
	NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_925__bF_buf0), .C(_526_), .Y(_855_) );
	NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1100__bF_buf1), .B(_855_), .C(_1551_), .Y(_856_) );
	MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(ABH_3_), .B(PC_11_), .S(_953__bF_buf4), .Y(_857_) );
	NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_928__bF_buf1), .B(_857_), .Y(_858_) );
	NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_858_), .C(_854_), .Y(_859_) );
	OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_674_), .C(_859_), .Y(_860_) );
	AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_850_), .C(_860_), .Y(_861_) );
	NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(PC_10_), .B(_670_), .C(_673_), .Y(_862_) );
	NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(PC_11_), .B(_670_), .C(_673_), .Y(_863_) );
	AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_862_), .C(_863_), .D(_859_), .Y(_864_) );
	INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_864_), .Y(_865_) );
	OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_840_), .C(RDY_bF_buf8), .Y(_866_) );
	OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_165_), .C(_866_), .D(_861_), .Y(_32_) );
	NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_840_), .Y(_867_) );
	NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_674_), .Y(_868_) );
	OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_1107_), .C(_1100__bF_buf0), .Y(_869_) );
	AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_1111_), .C(_869_), .Y(_870_) );
	NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_953__bF_buf3), .Y(_871_) );
	NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_939__bF_buf1), .Y(_872_) );
	OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_871_), .B(_872_), .C(_1479_), .Y(_873_) );
	AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_870_), .B(_873_), .Y(_874_) );
	OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_670_), .C(_874_), .Y(_875_) );
	OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_868_), .Y(_876_) );
	NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_867_), .Y(_877_) );
	NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_864_), .C(_818_), .Y(_878_) );
	INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_879_) );
	OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_878_), .C(RDY_bF_buf6), .Y(_880_) );
	OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_174_), .C(_880_), .D(_877_), .Y(_33_) );
	NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_695_), .Y(_881_) );
	OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_881_), .C(PC_13_), .Y(_882_) );
	OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(DIMUX_5_), .Y(_883_) );
	INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .Y(_884_) );
	AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ABH_5_), .C(_1237_), .Y(_885_) );
	OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_884_), .C(_885_), .Y(_886_) );
	AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(ABH_5_), .B(_708_), .C(_886_), .Y(_887_) );
	NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_887_), .C(_882_), .Y(_888_) );
	AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_876_), .C(_888_), .Y(_889_) );
	OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_875_), .C(_888_), .Y(_890_) );
	OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_890_), .B(_878_), .C(RDY_bF_buf4), .Y(_891_) );
	OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_178_), .C(_891_), .D(_889_), .Y(_34_) );
	NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_864_), .Y(_892_) );
	NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_892_), .C(_752_), .Y(_893_) );
	INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_894_) );
	OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_881_), .C(PC_14_), .Y(_895_) );
	INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_708_), .Y(_896_) );
	OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_1107_), .C(_1100__bF_buf3), .Y(_897_) );
	AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_1111_), .C(_897_), .Y(_898_) );
	OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_896_), .C(_898_), .Y(_899_) );
	AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_6_), .B(_676_), .C(_899_), .Y(_900_) );
	AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_900_), .C(_894_), .D(_893_), .Y(_901_) );
	AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_864_), .Y(_902_) );
	NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_902_), .C(_762_), .Y(_903_) );
	NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_900_), .Y(_904_) );
	NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_890_), .B(_904_), .C(_903_), .Y(_905_) );
	OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_905_), .C(RDY_bF_buf2), .Y(_906_) );
	OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_185_), .C(_906_), .Y(_35_) );
	NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_890_), .C(_840_), .Y(_907_) );
	NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_896_), .Y(_908_) );
	OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_881_), .C(PC_15_), .Y(_909_) );
	OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(DIMUX_7_), .Y(_910_) );
	OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_1107_), .C(_1100__bF_buf2), .Y(_911_) );
	AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_1111_), .C(_911_), .Y(_912_) );
	NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_912_), .C(_909_), .Y(_913_) );
	NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_908_), .B(_913_), .Y(_914_) );
	NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_914_), .C(_907_), .Y(_915_) );
	INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_916_) );
	NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_904_), .C(_893_), .Y(_917_) );
	AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_916_), .C(_924__bF_buf2), .Y(_918_) );
	AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(_190_), .C(_915_), .D(_918_), .Y(_36_) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .Y(AB_0_) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_1586_), .Y(AB_1_) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(AB_2_) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_1588_), .Y(AB_3_) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .Y(AB_4_) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .Y(AB_5_) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_1591_), .Y(AB_6_) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .Y(AB_7_) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .Y(AB_8_) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .Y(AB_9_) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .Y(AB_10_) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .Y(AB_11_) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(AB_12_) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .Y(AB_13_) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1584_), .Y(AB_14_) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .Y(AB_15_) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .Y(DO_0_) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .Y(DO_1_) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .Y(DO_2_) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .Y(DO_3_) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .Y(DO_4_) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(DO_5_) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .Y(DO_6_) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .Y(DO_7_) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(WE) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1371_), .Q(AXYS_0__0_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1388_), .Q(AXYS_0__1_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1395_), .Q(AXYS_0__2_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1402_), .Q(AXYS_0__3_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1406_), .Q(AXYS_0__4_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1418_), .Q(AXYS_0__5_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1424_), .Q(AXYS_0__6_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1432_), .Q(AXYS_0__7_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_111_), .Q(AXYS_1__0_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_114_), .Q(AXYS_1__1_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_117_), .Q(AXYS_1__2_) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_119_), .Q(AXYS_1__3_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_122_), .Q(AXYS_1__4_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_125_), .Q(AXYS_1__5_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_127_), .Q(AXYS_1__6_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_129_), .Q(AXYS_1__7_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_196_), .Q(AXYS_3__0_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_197_), .Q(AXYS_3__1_) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_199_), .Q(AXYS_3__2_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_202_), .Q(AXYS_3__3_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_205_), .Q(AXYS_3__4_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_208_), .Q(AXYS_3__5_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_211_), .Q(AXYS_3__6_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_214_), .Q(AXYS_3__7_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1553_), .Q(AXYS_2__0_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1556_), .Q(AXYS_2__1_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1559_), .Q(AXYS_2__2_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1562_), .Q(AXYS_2__3_) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1565_), .Q(AXYS_2__4_) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1567_), .Q(AXYS_2__5_) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1570_), .Q(AXYS_2__6_) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1573_), .Q(AXYS_2__7_) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_28_), .Q(NMI_edge) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(NMI), .Q(NMI_1) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_58_), .Q(cond_code_0_) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_59_), .Q(cond_code_1_) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_60_), .Q(cond_code_2_) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_72_), .Q(plp) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_71_), .Q(php) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_53_), .Q(clc) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_75_), .Q(sec) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_54_), .Q(cld) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_76_), .Q(sed) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_55_), .Q(cli) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_77_), .Q(sei) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_56_), .Q(clv) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_52_), .Q(bit_ins) );
	DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_67_), .Q(op_0_) );
	DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_68_), .Q(op_1_) );
	DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_69_), .Q(op_2_) );
	DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_70_), .Q(op_3_) );
	DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_74_), .Q(rotate) );
	DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_79_), .Q(shift_right) );
	DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_57_), .Q(compare) );
	DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_78_), .Q(shift) );
	DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_48_), .Q(adc_bcd) );
	DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_49_), .Q(adc_sbc) );
	DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_63_), .Q(inc) );
	DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_65_), .Q(load_only) );
	DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_83_), .Q(write_back) );
	DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_82_), .Q(store) );
	DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_64_), .Q(index_y) );
	DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_80_), .Q(src_reg_0_) );
	DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_81_), .Q(src_reg_1_) );
	DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_61_), .Q(dst_reg_0_) );
	DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_62_), .Q(dst_reg_1_) );
	DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_66_), .Q(load_reg) );
	DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_73_), .Q(res) );
	DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(DIMUX_0_), .Q(DIHOLD_0_) );
	DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(DIMUX_1_), .Q(DIHOLD_1_) );
	DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(DIMUX_2_), .Q(DIHOLD_2_) );
	DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(DIMUX_3_), .Q(DIHOLD_3_) );
	DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(DIMUX_4_), .Q(DIHOLD_4_) );
	DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(DIMUX_5_), .Q(DIHOLD_5_) );
	DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(DIMUX_6_), .Q(DIHOLD_6_) );
	DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(DIMUX_7_), .Q(DIHOLD_7_) );
	DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_18_), .Q(IRHOLD_0_) );
	DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_19_), .Q(IRHOLD_1_) );
	DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_20_), .Q(IRHOLD_2_) );
	DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_21_), .Q(IRHOLD_3_) );
	DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_22_), .Q(IRHOLD_4_) );
	DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_23_), .Q(IRHOLD_5_) );
	DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_24_), .Q(IRHOLD_6_) );
	DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_25_), .Q(IRHOLD_7_) );
	DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_26_), .Q(IRHOLD_valid) );
	DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_46_), .Q(V) );
	DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17_), .Q(D) );
	DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_27_), .Q(I) );
	DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_29_), .Q(N) );
	DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_47_), .Q(Z) );
	DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_16_), .Q(C) );
	DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_51_), .Q(backwards) );
	DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_50_), .Q(adj_bcd) );
	DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_8_), .Q(ABL_0_) );
	DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_9_), .Q(ABL_1_) );
	DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10_), .Q(ABL_2_) );
	DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_11_), .Q(ABL_3_) );
	DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_12_), .Q(ABL_4_) );
	DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_13_), .Q(ABL_5_) );
	DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_14_), .Q(ABL_6_) );
	DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_15_), .Q(ABL_7_) );
	DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0_), .Q(ABH_0_) );
	DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1_), .Q(ABH_1_) );
	DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2_), .Q(ABH_2_) );
	DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3_), .Q(ABH_3_) );
	DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4_), .Q(ABH_4_) );
	DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_5_), .Q(ABH_5_) );
	DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6_), .Q(ABH_6_) );
	DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_7_), .Q(ABH_7_) );
	DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_30_), .Q(PC_0_) );
	DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_37_), .Q(PC_1_) );
	DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_38_), .Q(PC_2_) );
	DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_39_), .Q(PC_3_) );
	DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_40_), .Q(PC_4_) );
	DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_41_), .Q(PC_5_) );
	DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_42_), .Q(PC_6_) );
	DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_43_), .Q(PC_7_) );
	DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_44_), .Q(PC_8_) );
	DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_45_), .Q(PC_9_) );
	DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_31_), .Q(PC_10_) );
	DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_32_), .Q(PC_11_) );
	DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_33_), .Q(PC_12_) );
	DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_34_), .Q(PC_13_) );
	DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_35_), .Q(PC_14_) );
	DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_36_), .Q(PC_15_) );
	DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_919_), .Q(state_0_), .R(_1257_), .S(vdd) );
	DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_920_), .Q(state_1_), .R(_1257_), .S(vdd) );
	DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_921_), .Q(state_2_), .R(_1257_), .S(vdd) );
	DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_922_), .Q(state_3_), .R(vdd), .S(_1257_) );
	DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_923_), .Q(state_4_), .R(_1257_), .S(vdd) );
	DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_931_), .Q(state_5_), .R(_1257_), .S(vdd) );
	OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(ADD_0_), .Y(_1783_) );
	NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(ADD_7_), .Y(_1784_) );
	NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(ADD_5_), .Y(_1785_) );
	NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(ADD_1_), .Y(_1786_) );
	NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1785_), .C(_1786_), .Y(_1787_) );
	NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1787_), .Y(ALU_Z) );
	INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(AI_7_), .Y(_1788_) );
	INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .Y(_1789_) );
	NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(ALU_AI7), .B(_1789__bF_buf3), .Y(_1790_) );
	OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1789__bF_buf2), .C(_1790_), .Y(_1604_) );
	NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(ALU_CI), .B(ALU_right), .Y(_1791_) );
	INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_1_), .Y(_1792_) );
	NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1792_), .Y(_1793_) );
	INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .Y(_1794_) );
	AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(ALU_BI_7_), .Y(_1795_) );
	NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(AI_7_), .B(_1795_), .Y(_1796_) );
	AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_7_), .B(_1792_), .C(_1793_), .D(_1796_), .Y(_1797_) );
	INVX4 INVX4_17 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .Y(_1798_) );
	OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(AI_7_), .B(_1795_), .C(_1798_), .Y(_1799_) );
	OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1797_), .C(_1791_), .Y(_1800_) );
	INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_2_), .Y(_1801_) );
	NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(_1801_), .Y(_1802_) );
	INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .Y(_1803_) );
	NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_7_), .B(_1803_), .Y(_1804_) );
	NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_op_2_), .Y(_1805_) );
	AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_7_), .B(_1805_), .C(_1804_), .Y(_1806_) );
	INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_1806_), .Y(_1807_) );
	INVX4 INVX4_18 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .Y(_1808_) );
	OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1806_), .Y(_1809_) );
	OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1807_), .C(_1809_), .Y(_1810_) );
	NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI7), .B(_1789__bF_buf1), .Y(_1811_) );
	OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf0), .B(_1810_), .C(_1811_), .Y(_1605_) );
	NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_1789__bF_buf3), .Y(_1812_) );
	OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(_1801_), .C(ALU_CI), .Y(_1813_) );
	NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(_1813_), .Y(_1814_) );
	NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_2_), .B(_1808_), .Y(_1815_) );
	NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_0_), .B(_1794_), .Y(_1816_) );
	NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_1_), .B(AI_0_), .Y(_1817_) );
	AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_0_), .B(_1817_), .C(_1793_), .D(_1816_), .Y(_1818_) );
	INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_0_), .Y(_1819_) );
	INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(AI_0_), .Y(_1820_) );
	OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1819_), .C(_1820_), .Y(_1821_) );
	NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1821_), .Y(_1822_) );
	NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(AI_1_), .Y(_1823_) );
	OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1822_), .C(_1823_), .Y(_1824_) );
	MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1805_), .S(_1819_), .Y(_1825_) );
	INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .Y(_1826_) );
	OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_1826_), .C(_1824_), .Y(_1617_) );
	MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_1_), .B(_1819_), .S(ALU_op_0_), .Y(_1618_) );
	NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_0_), .B(_1817_), .Y(_1619_) );
	NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(_1618_), .Y(_1620_) );
	AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1820_), .C(ALU_right), .Y(_1621_) );
	NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1620_), .Y(_1622_) );
	NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1825_), .C(_1622_), .Y(_1623_) );
	AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_1623_), .C(_1814_), .Y(_1624_) );
	INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .Y(_1625_) );
	OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1824_), .B(_1826_), .C(_1617_), .Y(_1626_) );
	OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1626_), .C(RDY_bF_buf8), .Y(_1627_) );
	OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1624_), .B(_1627_), .C(_1812_), .Y(_1609_) );
	NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_1789__bF_buf2), .Y(_1628_) );
	NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1824_), .Y(_1629_) );
	OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1629_), .C(_1617_), .Y(_1630_) );
	NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_1_), .B(_1794_), .Y(_1631_) );
	AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(ALU_BI_1_), .Y(_1632_) );
	INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(AI_1_), .Y(_1633_) );
	OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1633_), .C(ALU_BI_1_), .Y(_1634_) );
	OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1632_), .C(_1634_), .Y(_1635_) );
	NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_1_), .B(_1794_), .Y(_1636_) );
	AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1633_), .C(ALU_right), .Y(_1637_) );
	AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(AI_2_), .C(_1637_), .D(_1635_), .Y(_1638_) );
	OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_BI_1_), .C(_1801_), .Y(_1639_) );
	OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_1_), .B(_1803_), .C(_1639_), .Y(_1640_) );
	OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1640_), .Y(_1641_) );
	MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(_1640_), .S(_1638_), .Y(_1642_) );
	NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1642_), .B(_1630_), .Y(_1643_) );
	OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1825_), .Y(_1644_) );
	AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1824_), .B(_1644_), .C(_1814_), .D(_1623_), .Y(_1645_) );
	INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(AI_2_), .Y(_1646_) );
	NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_1_), .B(AI_1_), .Y(_1647_) );
	AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_1_), .B(_1647_), .C(_1793_), .D(_1636_), .Y(_1648_) );
	INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .Y(_1649_) );
	OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1646_), .C(_1648_), .D(_1649_), .Y(_1650_) );
	AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1640_), .Y(_1651_) );
	INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .Y(_1652_) );
	AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1640_), .C(_1650_), .Y(_1653_) );
	OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1651_), .C(_1645_), .Y(_1654_) );
	NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1654_), .Y(_1655_) );
	OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf1), .B(_1655_), .C(_1628_), .Y(_1610_) );
	NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_1789__bF_buf0), .Y(_1656_) );
	NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1640_), .B(_1650_), .Y(_1657_) );
	OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1645_), .C(_1657_), .Y(_1658_) );
	INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(AI_3_), .Y(_1659_) );
	INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_2_), .Y(_1660_) );
	NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1660_), .Y(_1661_) );
	OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1646_), .C(ALU_BI_2_), .Y(_1662_) );
	OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1661_), .C(_1662_), .Y(_1663_) );
	OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1660_), .C(_1646_), .Y(_1664_) );
	NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1664_), .C(_1663_), .Y(_1665_) );
	OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1659_), .C(_1665_), .Y(_1666_) );
	OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_BI_2_), .C(_1801_), .Y(_1667_) );
	OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_2_), .B(_1803_), .C(_1667_), .Y(_1668_) );
	NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1666_), .Y(_1669_) );
	NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(AI_3_), .Y(_1670_) );
	OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1668_), .Y(_1671_) );
	NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1670_), .B(_1665_), .C(_1671_), .Y(_1672_) );
	AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1672_), .Y(_1673_) );
	NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1673_), .B(_1658_), .Y(_1674_) );
	NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .B(_1669_), .Y(_1675_) );
	NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1675_), .C(_1643_), .Y(_1676_) );
	NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1676_), .Y(_1677_) );
	OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf3), .B(_1677_), .C(_1656_), .Y(_1611_) );
	NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_1789__bF_buf2), .Y(_1678_) );
	AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1668_), .C(_1673_), .D(_1658_), .Y(_1679_) );
	INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(AI_4_), .Y(_1680_) );
	INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_3_), .Y(_1681_) );
	NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1681_), .Y(_1682_) );
	OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1659_), .C(ALU_BI_3_), .Y(_1683_) );
	OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1682_), .C(_1683_), .Y(_1684_) );
	OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_0_), .B(_1681_), .C(_1659_), .Y(_1685_) );
	NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1685_), .C(_1684_), .Y(_1686_) );
	OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1680_), .C(_1686_), .Y(_1687_) );
	OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_BI_3_), .C(_1801_), .Y(_1688_) );
	OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_3_), .B(_1803_), .C(_1688_), .Y(_1689_) );
	NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1687_), .Y(_1690_) );
	AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1652_), .Y(_1691_) );
	OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1691_), .C(_1690_), .Y(_1692_) );
	XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(_1692_), .Y(_1693_) );
	OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf1), .B(_1693_), .C(_1678_), .Y(_1612_) );
	NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_1789__bF_buf0), .Y(_1694_) );
	NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1673_), .C(_1643_), .Y(_1695_) );
	NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .B(_1658_), .Y(_1696_) );
	NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1696_), .B(_1655_), .C(_1695_), .Y(_1697_) );
	NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(ALU_BCD), .B(_1697_), .Y(_1698_) );
	NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .B(_1679_), .Y(_1699_) );
	OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1691_), .C(_1699_), .Y(_1700_) );
	OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1693_), .C(_1700_), .Y(_1701_) );
	NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(AI_5_), .Y(_1702_) );
	AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(ALU_BI_4_), .Y(_1703_) );
	NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(AI_4_), .B(_1703_), .Y(_1704_) );
	AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(ALU_BI_4_), .C(_1793_), .D(_1704_), .Y(_1705_) );
	OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(AI_4_), .B(_1703_), .C(_1798_), .Y(_1706_) );
	OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1705_), .C(_1702_), .Y(_1707_) );
	NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_4_), .B(_1805_), .Y(_1708_) );
	OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_4_), .B(_1803_), .C(_1708_), .Y(_1709_) );
	OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_1709_), .C(_1707_), .Y(_1710_) );
	OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_1709_), .C(_1710_), .Y(_1711_) );
	INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .Y(_1712_) );
	NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1712_), .B(_1701_), .Y(_1713_) );
	OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1691_), .Y(_1714_) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(_1692_), .Y(_1715_) );
	INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(ALU_BCD), .Y(_1716_) );
	AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1677_), .B(_1655_), .C(_1716_), .Y(_1717_) );
	AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1699_), .C(_1715_), .D(_1717_), .Y(_1718_) );
	OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1718_), .C(RDY_bF_buf7), .Y(_1719_) );
	OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_1719_), .C(_1694_), .Y(_1613_) );
	NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .B(_1789__bF_buf3), .Y(_1720_) );
	OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1718_), .C(_1710_), .Y(_1721_) );
	NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(ALU_right), .B(AI_6_), .Y(_1722_) );
	AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(ALU_BI_5_), .Y(_1723_) );
	NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(AI_5_), .B(_1723_), .Y(_1724_) );
	AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(ALU_BI_5_), .C(_1793_), .D(_1724_), .Y(_1725_) );
	OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(AI_5_), .B(_1723_), .C(_1798_), .Y(_1726_) );
	OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1726_), .B(_1725_), .C(_1722_), .Y(_1727_) );
	OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_BI_5_), .C(_1801_), .Y(_1728_) );
	OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_5_), .B(_1803_), .C(_1728_), .Y(_1729_) );
	NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1727_), .Y(_1730_) );
	OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1729_), .Y(_1731_) );
	INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(_1731_), .Y(_1732_) );
	OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1732_), .C(_1730_), .Y(_1733_) );
	INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .Y(_1734_) );
	NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_1721_), .Y(_1735_) );
	INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .Y(_1736_) );
	OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(ALU_op_2_), .C(_1736_), .Y(_1737_) );
	AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_1737_), .C(_1712_), .D(_1701_), .Y(_1738_) );
	NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1738_), .Y(_1739_) );
	NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1735_), .Y(_1740_) );
	OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf2), .B(_1740_), .C(_1720_), .Y(_1614_) );
	NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_1789__bF_buf1), .Y(_1741_) );
	OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1738_), .C(_1730_), .Y(_1742_) );
	AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(ALU_BI_6_), .Y(_1743_) );
	NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(AI_6_), .B(_1743_), .Y(_1744_) );
	AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(ALU_BI_6_), .C(_1793_), .D(_1744_), .Y(_1745_) );
	OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(AI_6_), .B(_1743_), .C(_1798_), .Y(_1746_) );
	OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1798_), .C(_1746_), .D(_1745_), .Y(_1747_) );
	INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .Y(_1748_) );
	OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(ALU_BI_6_), .C(ALU_op_2_), .Y(_1749_) );
	OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI_6_), .B(_1748_), .C(_1749_), .Y(_1750_) );
	INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .Y(_1751_) );
	NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_1747_), .Y(_1752_) );
	NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(ALU_op_3_), .B(_1750_), .Y(_1753_) );
	OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_1753_), .C(_1752_), .Y(_1754_) );
	INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .Y(_1755_) );
	NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1742_), .Y(_1756_) );
	NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1754_), .C(_1735_), .Y(_1757_) );
	NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(_1756_), .Y(_1758_) );
	OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf0), .B(_1758_), .C(_1741_), .Y(_1615_) );
	INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .Y(_1759_) );
	AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1729_), .C(_1734_), .D(_1721_), .Y(_1760_) );
	OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .B(_1760_), .C(_1752_), .Y(_1761_) );
	OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_1807_), .C(_1800_), .Y(_1762_) );
	OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1807_), .C(_1762_), .Y(_1763_) );
	NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_1761_), .Y(_1764_) );
	INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .Y(_1765_) );
	NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1765_), .C(_1756_), .Y(_1766_) );
	NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1766_), .B(_1764_), .Y(_1767_) );
	NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1767_), .Y(_1768_) );
	OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .B(RDY_bF_buf5), .C(_1768_), .Y(_1616_) );
	NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(ALU_HC), .B(_1789__bF_buf3), .Y(_1769_) );
	OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf2), .B(_1718_), .C(_1769_), .Y(_1607_) );
	INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(ALU_N), .Y(_1770_) );
	OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1770_), .C(_1768_), .Y(_1608_) );
	NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1820_), .Y(_1771_) );
	INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .Y(_1772_) );
	AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1809_), .C(_1772_), .D(_1765_), .Y(_1773_) );
	NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1765_), .Y(_1774_) );
	OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1760_), .C(_1773_), .Y(_1775_) );
	NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_1775_), .Y(_1776_) );
	OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_1775_), .B(_1771_), .Y(_1777_) );
	AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1740_), .C(_1716_), .Y(_1778_) );
	AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1776_), .B(_1777_), .C(_1767_), .D(_1778_), .Y(_1779_) );
	NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(ALU_CO), .B(_1789__bF_buf1), .Y(_1780_) );
	OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1789__bF_buf0), .B(_1779_), .C(_1780_), .Y(_1606_) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ALU_AI7), .B(ALU_BI7), .Y(_1781_) );
	XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ALU_N), .B(ALU_CO), .Y(_1782_) );
	XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1781_), .B(_1782_), .Y(ALU_V) );
	DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1606_), .Q(ALU_CO) );
	DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1608_), .Q(ALU_N) );
	DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1607_), .Q(ALU_HC) );
	DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1609_), .Q(ADD_0_) );
	DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1610_), .Q(ADD_1_) );
	DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1611_), .Q(ADD_2_) );
	DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1612_), .Q(ADD_3_) );
	DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1613_), .Q(ADD_4_) );
	DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1614_), .Q(ADD_5_) );
	DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1615_), .Q(ADD_6_) );
	DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1616_), .Q(ADD_7_) );
	DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1605_), .Q(ALU_BI7) );
	DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1604_), .Q(ALU_AI7) );
endmodule
