module cpu ( gnd, vdd, clk, reset, DI, IRQ, NMI, RDY, AB, DO, WE);

input gnd, vdd;
input clk;
input reset;
input IRQ;
input NMI;
input RDY;
output WE;
input [7:0] DI;
output [15:0] AB;
output [7:0] DO;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf8) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf7) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf6) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf5) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf4) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf3) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf2) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf1) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(RDY), .Y(RDY_bF_buf0) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_799__bF_buf4) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_799__bF_buf3) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_799__bF_buf2) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_799__bF_buf1) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_799__bF_buf0) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf11) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf10) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf9) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf8) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1101__bF_buf3) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1101__bF_buf2) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1101__bF_buf1) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1101__bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_849_), .Y(_849__bF_buf4) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_849_), .Y(_849__bF_buf3) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_849_), .Y(_849__bF_buf2) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_849_), .Y(_849__bF_buf1) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_849_), .Y(_849__bF_buf0) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_825_), .Y(_825__bF_buf4) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_825_), .Y(_825__bF_buf3) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_825_), .Y(_825__bF_buf2) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_825_), .Y(_825__bF_buf1) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_825_), .Y(_825__bF_buf0) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf3) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf2) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf1) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf0) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_822_), .Y(_822__bF_buf4) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_822_), .Y(_822__bF_buf3) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_822_), .Y(_822__bF_buf2) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_822_), .Y(_822__bF_buf1) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_822_), .Y(_822__bF_buf0) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_152__bF_buf3) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_152__bF_buf2) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_152__bF_buf1) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_152__bF_buf0) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_795_), .Y(_795__bF_buf4) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_795_), .Y(_795__bF_buf3) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_795_), .Y(_795__bF_buf2) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_795_), .Y(_795__bF_buf1) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_795_), .Y(_795__bF_buf0) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_651_), .Y(_651__bF_buf4) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_651_), .Y(_651__bF_buf3) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_651_), .Y(_651__bF_buf2) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_651_), .Y(_651__bF_buf1) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_651_), .Y(_651__bF_buf0) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf4) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf3) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf2) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf1) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf0) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_830_), .Y(_830__bF_buf3) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_830_), .Y(_830__bF_buf2) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_830_), .Y(_830__bF_buf1) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_830_), .Y(_830__bF_buf0) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf3) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf2) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf1) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf0) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf7) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf6) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf5) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf4) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf3) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf2) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf1) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf0) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_859_), .Y(_859__bF_buf3) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_859_), .Y(_859__bF_buf2) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_859_), .Y(_859__bF_buf1) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_859_), .Y(_859__bF_buf0) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_148__bF_buf3) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_148__bF_buf2) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_148__bF_buf1) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_148__bF_buf0) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_815_), .Y(_815__bF_buf3) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_815_), .Y(_815__bF_buf2) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_815_), .Y(_815__bF_buf1) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_815_), .Y(_815__bF_buf0) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_812_), .Y(_812__bF_buf3) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_812_), .Y(_812__bF_buf2) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_812_), .Y(_812__bF_buf1) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_812_), .Y(_812__bF_buf0) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_809__bF_buf4) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_809__bF_buf3) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_809__bF_buf2) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_809__bF_buf1) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_809__bF_buf0) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(PC_13_), .Y(_787_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_788_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_789_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_790_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_790_), .Y(_791_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_791_), .Y(_792_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(_793_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_793_), .Y(_794_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(_794_), .Y(_795_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_792_), .Y(_796_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .Y(_797_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_797_), .Y(_798_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_798_), .Y(_799_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_800_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_800_), .Y(_801_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_802_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_801_), .Y(_803_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(_804_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_804_), .Y(_805_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_805_), .Y(_806_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf3), .B(_799__bF_buf4), .C(_803_), .D(_806_), .Y(_807_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_807_), .Y(_808_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(state_4_), .Y(_809_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_1_), .Y(_810_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_802_), .Y(_811_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(state_4_), .Y(_812_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_813_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_813_), .Y(_814_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf3), .B(_791_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf4), .B(_811_), .C(_815__bF_buf3), .Y(_816_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf2), .B(_805_), .C(_814_), .Y(_817_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf3), .B(_792_), .C(_817_), .Y(_818_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_818_), .Y(_819_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_819_), .Y(_820_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_820_), .Y(_821_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf1), .B(_810_), .C(_802_), .Y(_822_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(IRQ), .Y(_823_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(NMI_edge), .Y(_824_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(I), .B(_823_), .C(_824_), .Y(_825_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf4), .B(_822__bF_buf4), .Y(_826_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_821_), .C(PC_13_), .Y(_827_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(I), .Y(_828_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_824_), .Y(_829_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(NMI_edge), .C(_829_), .Y(_830_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_822__bF_buf3), .B(_830__bF_buf3), .Y(_831_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ABH_5_), .B(_831_), .Y(_832_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_804_), .Y(_833_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_833_), .Y(_834_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_834_), .Y(_835_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_813_), .Y(_836_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_837_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_836_), .Y(_838_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_798_), .C(_838_), .Y(_839_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_790_), .Y(_840_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_840_), .Y(_841_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_798_), .C(_841_), .Y(_842_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_839_), .C(_842_), .Y(_843_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_5_), .Y(_844_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(DI[5]), .Y(_845_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_844_), .C(_845_), .Y(DIMUX_5_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .Y(_846_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf0), .B(_789_), .C(_791_), .Y(_847_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_800_), .Y(_848_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf2), .B(_833_), .C(_848_), .Y(_849_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf1), .B(_840_), .C(_848_), .Y(_850_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf4), .B(ABH_5_), .C(_850_), .Y(_851_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_847_), .C(_851_), .Y(_852_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_5_), .C(_852_), .Y(_853_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_853_), .C(_827_), .Y(_854_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_808_), .C(_819_), .Y(_855_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_848_), .Y(_856_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf3), .B(_856_), .C(ADD_5_), .D(_849__bF_buf3), .Y(_857_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_812__bF_buf2), .C(_834_), .Y(_858_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(_822__bF_buf2), .Y(_859_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .Y(_860_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_825__bF_buf3), .Y(_861_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(ABL_5_), .Y(_862_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(IRQ), .B(_828_), .Y(_863_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_862_), .Y(_864_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_861_), .C(_859__bF_buf3), .Y(_865_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_865_), .C(_857_), .Y(_866_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .B(_843_), .C(_866_), .Y(_867_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_808_), .C(_819_), .Y(_868_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf2), .B(ADD_4_), .C(_850_), .Y(_869_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_847_), .Y(_870_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .B(_870_), .Y(_871_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(PC_4_), .Y(_872_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_825__bF_buf2), .Y(_873_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(ABL_4_), .Y(_874_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_874_), .Y(_875_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_873_), .C(_859__bF_buf2), .Y(_876_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_871_), .C(_869_), .Y(_877_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_843_), .C(_877_), .Y(_878_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_855_), .C(_868_), .D(_878_), .Y(_879_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .B(_808_), .C(_819_), .Y(_880_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf1), .B(_856_), .C(ADD_7_), .D(_849__bF_buf1), .Y(_881_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .B(_812__bF_buf0), .C(_834_), .Y(_882_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(PC_7_), .Y(_883_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_825__bF_buf1), .Y(_884_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(ABL_7_), .Y(_885_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_885_), .Y(_886_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_884_), .C(_859__bF_buf1), .Y(_887_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_887_), .C(_881_), .Y(_888_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_843_), .C(_888_), .Y(_889_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .B(_808_), .C(_819_), .Y(_890_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf0), .B(ADD_6_), .C(_850_), .Y(_891_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .B(_870_), .Y(_892_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(PC_6_), .Y(_893_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_825__bF_buf0), .Y(_894_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(ABL_6_), .Y(_895_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_895_), .Y(_896_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_894_), .C(_859__bF_buf0), .Y(_897_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_897_), .B(_892_), .C(_891_), .Y(_898_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_843_), .C(_898_), .Y(_899_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_889_), .B(_880_), .C(_890_), .D(_899_), .Y(_900_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_900_), .Y(_901_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(PC_0_), .B(_808_), .C(_819_), .Y(_902_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_807_), .C(ADD_0_), .Y(_903_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .Y(_904_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(PC_0_), .Y(_905_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_847_), .C(_904_), .D(_815__bF_buf2), .Y(_906_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(ABL_0_), .B(_825__bF_buf4), .Y(_907_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_825__bF_buf3), .C(_907_), .Y(_908_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf3), .B(_908_), .C(_906_), .Y(_909_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_903_), .Y(_910_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_842_), .Y(_911_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(CO), .B(backwards), .Y(_912_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_822__bF_buf1), .B(_825__bF_buf2), .C(_912_), .D(_815__bF_buf1), .Y(_913_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_3_), .Y(_914_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_814_), .Y(_915_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_812__bF_buf3), .C(_805_), .Y(_916_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf0), .B(_915_), .C(_916_), .Y(_917_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_913_), .C(_911_), .Y(_918_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_838_), .Y(_919_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_836_), .Y(_920_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_921_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf4), .B(_921_), .C(_919_), .Y(_922_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_914_), .Y(_923_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_923_), .Y(_924_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(_924_), .C(_812__bF_buf2), .Y(_925_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_792_), .C(_925_), .Y(_926_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_926_), .Y(_927_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_927_), .C(_902_), .D(_910_), .Y(_928_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_807_), .C(ADD_1_), .Y(_929_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(PC_1_), .B(_808_), .C(_819_), .Y(_930_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .Y(_931_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_815__bF_buf0), .C(res), .D(_817_), .Y(_932_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(PC_1_), .Y(_933_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_847_), .Y(_934_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_932_), .Y(_935_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(ABL_1_), .B(_825__bF_buf1), .Y(_936_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_825__bF_buf0), .C(_936_), .Y(_937_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf2), .B(_937_), .Y(_938_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_938_), .Y(_939_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_930_), .C(_939_), .Y(_940_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_808_), .C(_819_), .Y(_941_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf4), .B(ADD_3_), .C(_850_), .Y(_942_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .B(_870_), .Y(_943_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(PC_3_), .Y(_944_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_825__bF_buf4), .Y(_945_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(ABL_3_), .Y(_946_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_946_), .Y(_947_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_945_), .C(_859__bF_buf1), .Y(_948_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_943_), .C(_942_), .Y(_949_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_843_), .C(_949_), .Y(_950_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_808_), .C(_819_), .Y(_951_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(res), .B(_824_), .Y(_952_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_952_), .Y(_953_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf3), .B(ADD_2_), .C(_850_), .D(_953_), .Y(_954_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .B(_870_), .Y(_955_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(PC_2_), .Y(_956_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_825__bF_buf3), .Y(_957_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(ABL_2_), .Y(_958_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_958_), .Y(_959_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_957_), .C(_859__bF_buf0), .Y(_960_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_960_), .C(_954_), .Y(_961_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_843_), .C(_961_), .Y(_962_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_941_), .C(_951_), .D(_962_), .Y(_963_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_928_), .C(_963_), .Y(_964_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(PC_11_), .B(_808_), .C(_819_), .Y(_965_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_3_), .Y(_966_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(DI[3]), .Y(_967_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_966_), .C(_967_), .Y(DIMUX_3_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_812__bF_buf1), .C(_834_), .Y(_968_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf2), .B(ABH_3_), .C(_850_), .Y(_969_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(ABH_3_), .Y(_970_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_970_), .Y(_971_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(PC_11_), .Y(_972_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_825__bF_buf2), .Y(_973_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_973_), .C(_859__bF_buf3), .Y(_974_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_974_), .C(_969_), .Y(_975_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_3_), .C(_975_), .Y(_976_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(PC_10_), .B(_808_), .C(_819_), .Y(_977_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(DI[2]), .B(DIHOLD_2_), .S(RDY_bF_buf4), .Y(_978_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_978_), .Y(DIMUX_2_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_870_), .Y(_979_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf1), .B(ABH_2_), .C(_850_), .Y(_980_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(ABH_2_), .Y(_981_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_981_), .Y(_982_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(PC_10_), .Y(_983_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_825__bF_buf1), .Y(_984_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_984_), .C(_859__bF_buf2), .Y(_985_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_979_), .C(_980_), .Y(_986_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_2_), .C(_986_), .Y(_987_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_965_), .C(_977_), .D(_987_), .Y(_988_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(PC_9_), .B(_808_), .C(_819_), .Y(_989_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_1_), .Y(_990_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(DI[1]), .Y(_991_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_990_), .C(_991_), .Y(DIMUX_1_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_812__bF_buf0), .C(_834_), .Y(_992_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf0), .B(ABH_1_), .C(_850_), .Y(_993_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(ABH_1_), .Y(_994_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_994_), .Y(_995_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(PC_9_), .Y(_996_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_825__bF_buf0), .Y(_997_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_997_), .C(_859__bF_buf1), .Y(_998_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_992_), .B(_998_), .C(_993_), .Y(_999_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_1_), .C(_999_), .Y(_1000_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .B(_808_), .C(_819_), .Y(_1001_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(DIHOLD_0_), .Y(_1002_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(DI[0]), .Y(_1003_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1002_), .C(_1003_), .Y(DIMUX_0_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_870_), .Y(_1004_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf4), .B(ABH_0_), .C(_850_), .Y(_1005_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(ABH_0_), .Y(_1006_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_824_), .C(_1006_), .Y(_1007_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .Y(_1008_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_825__bF_buf4), .Y(_1009_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_1009_), .C(_859__bF_buf0), .Y(_1010_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1004_), .C(_1005_), .Y(_1011_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_0_), .C(_1011_), .Y(_1012_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_989_), .C(_1001_), .D(_1012_), .Y(_1013_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_1013_), .Y(_1014_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_1014_), .C(_964_), .Y(_1015_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(PC_12_), .Y(_1016_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .Y(_1017_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(DIHOLD_4_), .Y(_1018_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf7), .B(DI[4]), .C(_1018_), .Y(_1019_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(DIMUX_4_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(ABH_4_), .Y(_1020_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_815__bF_buf3), .C(_817_), .Y(_1021_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_870_), .C(_1021_), .Y(_1022_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_825__bF_buf3), .Y(_1023_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_830__bF_buf2), .Y(_1024_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1024_), .C(_859__bF_buf3), .Y(_1025_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1022_), .Y(_1026_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(DIMUX_4_), .C(_1026_), .Y(_1027_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_820_), .C(_1027_), .Y(_1028_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1028_), .C(_854_), .Y(_1029_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_900_), .Y(_1030_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_928_), .Y(_1031_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_941_), .Y(_1032_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_807_), .C(ADD_3_), .Y(_1033_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_943_), .Y(_1034_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_948_), .C(_1034_), .Y(_1035_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_951_), .Y(_1036_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_807_), .C(ADD_2_), .Y(_1037_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_955_), .Y(_1038_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_960_), .C(_1038_), .Y(_1039_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1032_), .C(_1036_), .D(_1039_), .Y(_1040_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .B(_1031_), .Y(_1041_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_1013_), .Y(_1042_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1042_), .C(_1041_), .Y(_1043_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_854_), .Y(_1044_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_1043_), .C(RDY_bF_buf6), .Y(_1045_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(RDY_bF_buf5), .C(_1029_), .D(_1045_), .Y(_9__13_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(PC_14_), .B(_1017__bF_buf6), .Y(_1046_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_1043_), .Y(_1047_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_821_), .C(PC_14_), .Y(_1048_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(ABH_6_), .Y(_1049_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_815__bF_buf2), .C(_817_), .Y(_1050_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_870_), .C(_1050_), .Y(_1051_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(DI[6]), .B(DIHOLD_6_), .S(RDY_bF_buf4), .Y(_1052_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1052_), .Y(DIMUX_6_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(ABH_6_), .B(_831_), .C(DIMUX_6_), .D(_843_), .Y(_1053_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1053_), .C(_1048_), .Y(_1054_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1047_), .Y(_1055_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_1028_), .Y(_1056_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1054_), .C(_1015_), .Y(_1057_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1057_), .Y(_1058_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1055_), .C(_1046_), .Y(_9__14_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(PC_15_), .Y(_1059_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_821_), .C(PC_15_), .Y(_1060_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(ABH_7_), .Y(_1061_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_815__bF_buf1), .C(_817_), .Y(_1062_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(ABH_7_), .B(_831_), .C(_1062_), .Y(_1063_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(DI[7]), .B(DIHOLD_7_), .S(RDY_bF_buf2), .Y(_1064_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .Y(DIMUX_7_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_870_), .C(DIMUX_7_), .D(_843_), .Y(_1065_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1065_), .C(_1060_), .Y(_1066_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1067_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1067_), .C(_1047_), .Y(_1068_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1066_), .C(_1017__bF_buf5), .Y(_1069_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf4), .B(_1059_), .C(_1068_), .D(_1069_), .Y(_9__15_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_822__bF_buf0), .Y(_1070_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_801_), .Y(_1071_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf3), .B(_1071_), .Y(_1072_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .Y(_1073_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_3_), .Y(_1074_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(DIMUX_3_), .Y(_1075_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1074_), .C(_1075_), .Y(_1076_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf1), .B(_1076_), .Y(_1077_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_2_), .Y(_1078_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_978_), .C(_1078_), .Y(_1079_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(_830__bF_buf0), .Y(_1080_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1077_), .Y(_1081_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .B(IRHOLD_1_), .S(_1073_), .Y(_1082_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf2), .B(_1082_), .Y(_1083_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(IRHOLD_0_), .S(_1073_), .Y(_1084_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf1), .B(_1084_), .Y(_1085_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1085_), .Y(_1086_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1086_), .B(_1081_), .Y(_1087_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_7_), .Y(_1088_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_1064_), .C(_1088_), .Y(_1089_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf3), .B(_1089_), .Y(_1090_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_4_), .Y(_1091_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_1019_), .C(_1091_), .Y(_1092_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .B(IRHOLD_5_), .S(_1073_), .Y(_1093_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf0), .B(_1093_), .Y(_1094_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf2), .B(_1092_), .C(_1094_), .Y(_1095_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1095_), .Y(_1096_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1087_), .Y(_1097_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1072_), .C(_1070__bF_buf4), .D(_1097_), .Y(_1098_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf3), .B(_921_), .Y(_1099_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .Y(_1100_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .Y(_1101_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_830__bF_buf1), .Y(_1102_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(_1076_), .C(_830__bF_buf0), .Y(_1103_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1103_), .C(_1086_), .Y(_1104_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1100_), .C(_1101__bF_buf3), .D(_1104_), .Y(_1105_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_1106_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_1106_), .Y(_1107_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_793_), .Y(_1108_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1107_), .Y(_1109_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_914_), .C(_1108_), .Y(_1110_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .Y(_1111_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1109_), .C(_1112_), .Y(_1113_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1107_), .Y(_1114_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_924_), .Y(_1115_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1115_), .S(_1017__bF_buf1), .Y(_1116_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_1113_), .Y(_1117_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_806_), .C(_1017__bF_buf0), .Y(_1118_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_805_), .Y(_1119_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf1), .B(_1119_), .C(RDY_bF_buf7), .Y(_1120_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1120_), .Y(_1121_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf3), .B(_841_), .Y(_1122_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf2), .B(_1119_), .Y(_1123_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1123_), .Y(_1124_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1122_), .C(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1125_), .Y(_1126_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf2), .B(_1119_), .Y(_1127_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf1), .B(_806_), .C(_1017__bF_buf7), .Y(_1128_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf6), .B(_1127_), .C(_1128_), .Y(_1129_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf1), .B(_1071_), .Y(_1130_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf0), .B(_923_), .C(RDY_bF_buf4), .Y(_1131_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1130_), .C(_1131_), .Y(_1132_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1132_), .Y(_1133_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1117_), .C(_1126_), .Y(_1134_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1134_), .B(_1105_), .Y(_1135_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_1076_), .C(_830__bF_buf3), .Y(_1136_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_837_), .Y(_1137_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .Y(_1138_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf0), .B(_1138_), .Y(_1139_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf2), .B(_1079_), .Y(_1140_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1101__bF_buf2), .Y(_1141_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_1139_), .C(_1136_), .D(_1141_), .Y(_1142_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf2), .B(_1137_), .Y(_1143_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1144_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_814_), .Y(_1145_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf4), .B(_1145_), .C(RDY_bF_buf2), .Y(_1146_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1144_), .C(_1146_), .Y(_1147_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1142_), .Y(_1148_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_848_), .Y(_1149_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1149_), .Y(_1150_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1150_), .Y(_1151_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_796_), .C(_1151_), .Y(_1152_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .Y(_1153_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_1149_), .Y(_1154_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf4), .B(_792_), .Y(_1155_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf4), .B(_1155_), .Y(_1156_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1154_), .C(_1156_), .Y(_1157_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1157_), .Y(_1158_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1158_), .Y(_1159_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_856_), .Y(_1160_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_805_), .Y(_1161_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf3), .B(_1161_), .Y(_1162_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1162_), .Y(_1163_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_1160_), .C(_1163_), .Y(_1164_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_916_), .S(RDY_bF_buf7), .Y(_1165_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1165_), .Y(_1166_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_912_), .Y(_1167_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_847_), .C(_815__bF_buf0), .D(_1167_), .Y(_1168_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .Y(_1169_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf0), .B(_1161_), .Y(_1170_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_814_), .Y(_1171_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_1171_), .C(RDY_bF_buf4), .Y(_1172_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1170_), .C(_1172_), .Y(_1173_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1169_), .Y(_1174_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_1166_), .Y(_1176_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1159_), .Y(_1177_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf1), .B(_1092_), .Y(_1178_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_3_), .Y(_1179_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(IRHOLD_3_), .C(_830__bF_buf0), .Y(_1180_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1179_), .C(_1180_), .Y(_1181_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1181_), .Y(_1182_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf4), .B(_1082_), .C(_1085_), .Y(_1183_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1182_), .Y(_1184_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1184_), .Y(_1185_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1077_), .Y(_1186_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1102_), .Y(_1187_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf3), .B(_1084_), .C(_1187_), .Y(_1188_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1188_), .C(_1185_), .Y(_1189_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_1107_), .C(_794_), .Y(_1190_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .Y(_1191_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_1191_), .Y(_1192_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_1190_), .C(_1192_), .Y(_1193_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf3), .B(_1071_), .C(_1109_), .Y(_1194_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_813_), .Y(_1195_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_1195_), .Y(_1196_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf1), .B(_1196_), .Y(_1197_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_1138_), .C(_1197_), .Y(_1198_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1194_), .Y(_1199_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_1193_), .C(_1199_), .Y(_1200_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_810_), .C(_798_), .Y(_1201_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .Y(_1202_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1202_), .Y(_1203_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_919_), .C(_1203_), .Y(_1204_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf0), .B(_838_), .Y(_1205_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1196_), .Y(_1206_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(store), .B(CO), .Y(_1207_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1207_), .Y(_1208_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1205_), .C(_1208_), .D(_1206_), .Y(_1209_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_1106_), .Y(_1210_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf3), .B(_1210_), .Y(_1211_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(write_back), .Y(_1212_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1212_), .Y(_1213_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1213_), .Y(_1214_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1211_), .Y(_1215_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1209_), .Y(_1216_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1216_), .Y(_1217_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(_1198_), .Y(_1218_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1212_), .C(_1218_), .Y(_1219_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1219_), .C(_1217_), .Y(_1220_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1070__bF_buf2), .C(_1220_), .Y(_1221_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1086_), .Y(_1222_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1092_), .C(_830__bF_buf3), .Y(_1223_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(IRHOLD_6_), .Y(_1224_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_1052_), .C(_1224_), .Y(_1225_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_830__bF_buf2), .B(_1225_), .Y(_1226_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1094_), .Y(_1227_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1227_), .Y(_1228_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf1), .B(_1228_), .C(_1222_), .Y(_1229_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_798_), .C(_801_), .Y(_1230_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1230_), .Y(_1231_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1206_), .C(RDY_bF_buf3), .Y(_1232_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf3), .B(_921_), .C(_1017__bF_buf0), .Y(_1233_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1233_), .Y(_1234_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_1234_), .C(_1229_), .Y(_1235_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_789_), .Y(_1236_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_799__bF_buf1), .Y(_1237_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf7), .B(_1237_), .Y(_1238_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(write_back), .C(_1218_), .Y(_1239_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_795__bF_buf2), .Y(_1240_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf1), .B(_915_), .C(RDY_bF_buf1), .Y(_1241_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1240_), .C(_1241_), .Y(_1242_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1242_), .C(_1239_), .Y(_1243_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_810_), .C(_794_), .Y(_1244_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .Y(_1245_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf0), .B(_803_), .C(_1017__bF_buf6), .Y(_1246_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_1245_), .C(_1246_), .Y(_1247_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf2), .B(_915_), .Y(_1248_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf1), .B(_1236_), .C(_1017__bF_buf4), .Y(_1249_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1248_), .C(_1249_), .Y(_1250_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_1145_), .Y(_1251_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf3), .B(_1138_), .C(_1017__bF_buf2), .Y(_1252_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_1251_), .C(_1252_), .Y(_1253_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1250_), .C(_1253_), .Y(_1254_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1243_), .Y(_1255_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(_1235_), .C(_1221_), .Y(_1256_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1256_), .Y(_1257_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1135_), .C(_1257_), .Y(_1438__0_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .Y(_1258_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1253_), .C(_1258_), .Y(_1259_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1259_), .Y(_1260_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1251_), .Y(_1261_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_0_), .Y(_1262_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(_1262_), .C(_825__bF_buf2), .Y(_1263_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_valid), .B(DIMUX_0_), .C(_1263_), .Y(_1264_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf1), .B(_1082_), .C(_1264_), .Y(_1265_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1182_), .Y(_1266_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_830__bF_buf1), .Y(_1267_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1178_), .Y(_1268_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1268_), .Y(_1269_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_1269_), .C(_1266_), .Y(_1270_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf0), .B(_1145_), .C(_1017__bF_buf7), .Y(_1271_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf6), .B(_1237_), .C(_1271_), .Y(_1272_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1272_), .C(_1270_), .Y(_1273_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1178_), .Y(_1274_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_830__bF_buf0), .Y(_1275_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf0), .B(_1093_), .C(_1275_), .Y(_1276_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1274_), .Y(_1277_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1181_), .Y(_1278_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1278_), .Y(_1279_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1277_), .Y(_1280_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf2), .B(_806_), .C(_916_), .Y(_1281_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1281_), .Y(_1282_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1150_), .C(_1282_), .Y(_1283_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1070__bF_buf0), .C(_1283_), .Y(_1284_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf0), .B(_1145_), .Y(_1285_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_1285_), .Y(_1286_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1186_), .Y(_1287_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(_1178_), .Y(_1288_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_1288_), .Y(_1289_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1289_), .C(_1284_), .Y(_1290_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf1), .B(_1171_), .Y(_1291_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1094_), .Y(_1292_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .Y(_1293_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1293_), .Y(_1294_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1294_), .Y(_1295_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf4), .B(_1291_), .C(_1070__bF_buf3), .D(_1295_), .Y(_1296_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .Y(_1297_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1186_), .Y(_1298_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1094_), .Y(_1299_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1274_), .Y(_1300_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1300_), .Y(_1301_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1297_), .C(_1070__bF_buf2), .D(_1301_), .Y(_1302_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(Z), .Y(_1303_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_1303_), .Y(_1304_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(C), .C(_1304_), .Y(_1305_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(V), .Y(_1306_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_1306_), .Y(_1307_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(N), .C(_1307_), .Y(_1308_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_1308_), .S(cond_code_2_), .Y(_1309_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(cond_code_0_), .Y(_1310_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1099_), .C(_1310_), .Y(_1311_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .Y(_1312_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1312_), .Y(_1313_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1154_), .C(_1313_), .Y(_1314_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_849__bF_buf3), .C(_1314_), .Y(_1315_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1315_), .Y(_1316_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1302_), .C(_1296_), .Y(_1317_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_1290_), .C(_1317_), .Y(_1318_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_915_), .Y(_1319_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1319_), .Y(_1320_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(RDY_bF_buf3), .Y(_1321_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1070__bF_buf1), .C(_1287_), .Y(_1322_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf4), .B(_915_), .Y(_1323_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf3), .B(_1071_), .C(RDY_bF_buf2), .Y(_1324_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_1323_), .C(_1324_), .Y(_1325_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_850_), .Y(_1326_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1122_), .C(_1326_), .Y(_1327_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf7), .B(_1248_), .C(_1327_), .Y(_1328_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1328_), .Y(_1329_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1182_), .C(_1278_), .Y(_1330_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf0), .B(_1178_), .Y(_1331_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(_1331_), .C(_1329_), .Y(_1332_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1322_), .C(_1332_), .Y(_1333_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .Y(_1334_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1334_), .C(_1318_), .Y(_1438__1_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf4), .B(_811_), .C(_1017__bF_buf6), .Y(_1335_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_792_), .Y(_1336_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_841_), .C(_1336_), .Y(_1337_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .Y(_1338_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1338_), .Y(_1339_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_924_), .C(_798_), .Y(_1340_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1337_), .C(_1339_), .Y(_1341_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_815__bF_buf3), .Y(_1342_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_1342_), .Y(_1343_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .B(_1310_), .C(_1343_), .Y(_1344_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_1341_), .Y(_1345_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1181_), .Y(_1346_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf3), .B(_1346_), .Y(_1347_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1087_), .C(_1347_), .Y(_1348_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1277_), .C(_1298_), .Y(_1349_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1274_), .Y(_1350_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1277_), .C(_1298_), .D(_1350_), .Y(_1351_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(_1178_), .C(_1298_), .D(_1300_), .Y(_1352_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_1351_), .C(_1352_), .Y(_1353_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1353_), .Y(_1354_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf4), .B(_1084_), .C(_1267_), .Y(_1355_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1355_), .Y(_1356_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1103_), .C(_1178_), .D(_1184_), .Y(_1357_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf3), .B(_1084_), .C(_1083_), .Y(_1358_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1182_), .Y(_1359_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1274_), .C(_1359_), .Y(_1360_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_825__bF_buf2), .Y(_1361_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1361_), .Y(_1362_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1265_), .C(_1182_), .Y(_1363_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1330_), .C(_1362_), .D(_1363_), .Y(_1364_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1360_), .C(_1364_), .Y(_1365_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1090_), .C(_1102_), .Y(_1366_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1183_), .Y(_1367_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1278_), .Y(_1368_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1366_), .C(_1367_), .D(_1368_), .Y(_1369_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1225_), .C(_830__bF_buf3), .Y(_1370_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1370_), .C(_1298_), .Y(_1371_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1300_), .C(_1102_), .D(_1287_), .Y(_1372_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .B(_1369_), .C(_1372_), .Y(_1373_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1365_), .Y(_1374_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1345_), .C(_1354_), .D(_1374_), .Y(_1375_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .Y(_1376_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf0), .B(_1376_), .C(_1017__bF_buf4), .Y(_1377_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1240_), .C(_1377_), .Y(_1378_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_1161_), .C(RDY_bF_buf0), .Y(_1380_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1245_), .C(_1380_), .Y(_1381_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_1161_), .C(RDY_bF_buf7), .Y(_1382_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1202_), .C(_1382_), .Y(_1383_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1383_), .B(_1381_), .Y(_1384_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1379_), .Y(_1385_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(_1385_), .Y(_1386_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1273_), .Y(_1387_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .Y(_1388_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1388_), .Y(_1389_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1087_), .C(_1389_), .Y(_1390_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_1390_), .Y(_1391_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf1), .B(_1376_), .Y(_1392_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1392_), .Y(_1393_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .Y(_1394_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_1211_), .C(RDY_bF_buf5), .Y(_1395_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_1394_), .C(_1395_), .Y(_1396_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1396_), .C(_1391_), .Y(_1397_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1253_), .C(_1169_), .Y(_1398_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1105_), .Y(_1399_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1159_), .C(_1399_), .Y(_1400_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1400_), .Y(_1401_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1235_), .C(_1401_), .Y(_1402_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1402_), .Y(_1403_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1403_), .Y(_1438__2_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .Y(_1404_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_1300_), .C(_1279_), .Y(_1405_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_1404_), .C(_1405_), .Y(_1406_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf0), .B(_1119_), .C(_1017__bF_buf1), .Y(_1407_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf4), .B(_792_), .C(RDY_bF_buf2), .Y(_1408_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1408_), .C(_1406_), .Y(_1409_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .Y(_1410_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1111_), .C(_1331_), .D(_1346_), .Y(_1411_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_795__bF_buf3), .C(_1017__bF_buf7), .Y(_1412_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf6), .B(_1144_), .C(_1412_), .Y(_1413_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(_1411_), .Y(_1414_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_812__bF_buf2), .B(_924_), .Y(_1415_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_799__bF_buf3), .Y(_1416_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf2), .B(_1138_), .C(RDY_bF_buf1), .Y(_1417_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_1416_), .C(_1417_), .Y(_1418_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_1415_), .C(_1418_), .Y(_1419_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_1414_), .Y(_1420_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf2), .B(_1369_), .C(_1420_), .Y(_1421_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1410_), .Y(_1422_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1135_), .Y(_1423_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1397_), .C(_1423_), .Y(_1424_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_1424_), .C(_1318_), .Y(_1425_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1375_), .C(_1257_), .Y(_1426_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1344_), .C(_1335_), .Y(_1427_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_1374_), .Y(_1428_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1428_), .Y(_1429_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1287_), .Y(_1430_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf1), .B(_1430_), .C(_1286_), .Y(_1431_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1253_), .Y(_1432_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1129_), .Y(_1433_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1432_), .Y(_1434_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(_1121_), .Y(_1435_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .B(_1435_), .Y(_1436_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1166_), .Y(_1437_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1437_), .C(_1436_), .Y(_41_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1431_), .C(_41_), .Y(_42_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .Y(_43_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1298_), .Y(_44_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_43_), .C(_1101__bF_buf0), .D(_44_), .Y(_45_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1298_), .Y(_46_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1160_), .C(_1101__bF_buf3), .D(_46_), .Y(_47_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_45_), .C(_47_), .Y(_48_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1409_), .Y(_49_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_48_), .C(_49_), .Y(_50_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_1429_), .Y(_51_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .B(_1426_), .C(_51_), .Y(_1438__3_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .Y(_52_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1152_), .C(_52_), .Y(_53_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_1381_), .Y(_54_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_54_), .C(_1434_), .Y(_55_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_53_), .Y(_56_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_56_), .Y(_57_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_1320_), .C(_1322_), .Y(_58_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_58_), .Y(_59_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1270_), .C(_1284_), .Y(_60_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_60_), .Y(_61_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_59_), .C(_61_), .Y(_1438__4_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_1238_), .Y(_62_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .Y(_63_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_63_), .Y(_64_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_65_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1113_), .Y(_67_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1157_), .Y(_68_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_67_), .Y(_69_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_66_), .C(_69_), .Y(_70_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .Y(_71_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1408_), .C(_71_), .Y(_72_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_1383_), .C(_72_), .Y(_73_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_70_), .Y(_74_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_1411_), .C(_74_), .Y(_75_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_1229_), .Y(_76_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1302_), .C(_76_), .Y(_77_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_75_), .Y(_78_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1393_), .C(_78_), .Y(_1438__5_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(C), .Y(_79_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_1210_), .C(_798_), .Y(_80_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_803_), .B(_809__bF_buf3), .C(_80_), .Y(_81_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(load_only), .Y(_82_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(shift), .B(_82_), .Y(_83_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(rotate), .B(_81_), .C(_83_), .Y(_84_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(rotate), .Y(_85_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(compare), .Y(_86_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(shift), .Y(_87_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_88_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(inc), .B(_87_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_1205_), .C(_89_), .Y(_90_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .Y(_91_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf2), .B(_1236_), .C(_815__bF_buf2), .Y(_92_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .C(CO), .Y(_93_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_1161_), .C(_1154_), .Y(_94_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf1), .B(_1171_), .C(_1230_), .Y(_95_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_95_), .Y(_96_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .Y(_97_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf0), .B(_792_), .C(_1143_), .Y(_98_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_99_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_97_), .C(_99_), .Y(_100_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_96_), .Y(_101_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_101_), .Y(_102_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_90_), .C(_102_), .Y(_103_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_84_), .C(_103_), .Y(CI) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .Y(_104_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_88_), .Y(_105_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_812__bF_buf1), .C(_1170_), .Y(_106_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf2), .B(_1245_), .Y(_107_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_106_), .Y(_108_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_1195_), .Y(_109_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_109_), .C(_812__bF_buf0), .Y(_110_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1251_), .Y(_111_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .Y(_112_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_112_), .Y(_113_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .Y(_114_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_99_), .C(_1100_), .Y(_115_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_115_), .Y(_116_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_113_), .C(_116_), .Y(_117_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_1100_), .C(_104_), .D(_117_), .Y(BI_0_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .Y(_118_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_1100_), .C(_118_), .D(_117_), .Y(BI_1_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_1100_), .C(_978_), .D(_117_), .Y(BI_2_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_1100_), .C(_1179_), .D(_117_), .Y(BI_3_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_1100_), .C(_1019_), .D(_117_), .Y(BI_4_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .Y(_119_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_1100_), .C(_119_), .D(_117_), .Y(BI_5_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_1100_), .C(_1052_), .D(_117_), .Y(BI_6_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_1100_), .C(_1064_), .D(_117_), .Y(BI_7_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_815__bF_buf1), .Y(_120_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf1), .B(_1171_), .C(_106_), .Y(_121_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_94_), .Y(_122_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_122_), .C(ADD_0_), .Y(_123_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf4), .B(_1236_), .C(_1100_), .Y(_124_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_125_), .C(_123_), .Y(_126_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_126_), .Y(_127_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(src_reg_1_), .Y(_128_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf0), .B(_915_), .C(_1110_), .Y(_129_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf1), .B(_1236_), .C(_809__bF_buf4), .D(_1145_), .Y(_130_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf2), .B(_129_), .C(_130_), .Y(_131_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf3), .B(_1119_), .C(_795__bF_buf0), .D(_1171_), .Y(_132_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf3), .B(_1119_), .C(_1160_), .Y(_133_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_133_), .Y(_134_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_1145_), .C(_916_), .Y(_135_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1137_), .Y(_136_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_915_), .C(_136_), .Y(_137_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1244_), .C(_1230_), .Y(_138_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_135_), .C(_138_), .Y(_139_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_139_), .C(_134_), .Y(_140_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_1_), .Y(_141_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .Y(_142_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_822__bF_buf4), .C(_142_), .Y(_143_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_140_), .C(_144_), .Y(_145_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__0_), .Y(_147_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(src_reg_0_), .Y(_148_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf2), .B(_811_), .C(_142_), .Y(_149_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .C(index_y), .Y(_150_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_0_), .B(_859__bF_buf1), .Y(_151_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .C(_149_), .Y(_152_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_152__bF_buf3), .C(_148__bF_buf3), .Y(_153_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__0_), .Y(_154_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(src_reg_0_), .B(_140_), .C(_152__bF_buf2), .Y(_155_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_155__bF_buf3), .Y(_156_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_156_), .C(_153_), .Y(_157_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__0_), .Y(_158_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_152__bF_buf1), .C(_148__bF_buf2), .Y(_159_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__0_), .Y(_160_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_155__bF_buf2), .Y(_161_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_161_), .C(_159_), .Y(_162_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_162_), .Y(_163_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1123_), .Y(_164_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_1319_), .C(_798_), .Y(_165_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_798_), .C(_856_), .Y(_166_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_164_), .C(_167_), .Y(_168_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .Y(_169_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_1251_), .Y(_170_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_142_), .Y(_171_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_168_), .Y(_172_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_163_), .C(_127_), .Y(AI_0_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_98_), .Y(_173_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_815__bF_buf0), .C(_118_), .D(_125_), .Y(_174_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_1_), .C(_174_), .Y(_175_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__1_), .Y(_176_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_177_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__1_), .Y(_178_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_155__bF_buf1), .Y(_179_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_179_), .C(_177_), .Y(_180_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__1_), .Y(_181_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_152__bF_buf3), .C(_148__bF_buf0), .Y(_182_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__1_), .Y(_183_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_155__bF_buf0), .Y(_184_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_184_), .C(_182_), .Y(_185_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_185_), .Y(_186_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_186_), .C(_175_), .Y(AI_1_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_815__bF_buf3), .C(_978_), .D(_125_), .Y(_187_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_2_), .C(_187_), .Y(_188_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__2_), .Y(_189_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_190_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__2_), .Y(_191_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_155__bF_buf3), .Y(_192_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_192_), .C(_190_), .Y(_193_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__2_), .Y(_194_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_152__bF_buf1), .C(_148__bF_buf2), .Y(_195_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__2_), .Y(_196_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_155__bF_buf2), .Y(_197_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_197_), .C(_195_), .Y(_198_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_198_), .Y(_199_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_199_), .C(_188_), .Y(AI_2_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_815__bF_buf2), .C(_1179_), .D(_125_), .Y(_200_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_3_), .C(_200_), .Y(_201_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__3_), .Y(_202_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_203_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__3_), .Y(_204_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_155__bF_buf1), .Y(_205_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_205_), .C(_203_), .Y(_206_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__3_), .Y(_207_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_152__bF_buf3), .C(_148__bF_buf0), .Y(_208_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__3_), .Y(_209_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_155__bF_buf0), .Y(_210_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_210_), .C(_208_), .Y(_211_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_211_), .Y(_212_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_212_), .C(_201_), .Y(AI_3_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_815__bF_buf1), .C(_1019_), .D(_125_), .Y(_213_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_4_), .C(_213_), .Y(_214_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__4_), .Y(_215_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_216_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__4_), .Y(_217_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_155__bF_buf3), .Y(_218_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_218_), .C(_216_), .Y(_219_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__4_), .Y(_220_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_152__bF_buf1), .C(_148__bF_buf2), .Y(_221_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__4_), .Y(_222_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_155__bF_buf2), .Y(_223_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_223_), .C(_221_), .Y(_224_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_224_), .Y(_225_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_225_), .C(_214_), .Y(AI_4_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(ABH_5_), .Y(_226_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_815__bF_buf0), .C(_119_), .D(_125_), .Y(_227_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_5_), .C(_227_), .Y(_228_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__5_), .Y(_229_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_230_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__5_), .Y(_231_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_155__bF_buf1), .Y(_232_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_232_), .C(_230_), .Y(_233_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__5_), .Y(_234_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_152__bF_buf3), .C(_148__bF_buf0), .Y(_235_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__5_), .Y(_236_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_155__bF_buf0), .Y(_237_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_237_), .C(_235_), .Y(_238_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_238_), .Y(_239_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_239_), .C(_228_), .Y(AI_5_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_815__bF_buf3), .C(_1052_), .D(_125_), .Y(_240_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_6_), .C(_240_), .Y(_241_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__6_), .Y(_242_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_243_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__6_), .Y(_244_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_155__bF_buf3), .Y(_245_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_245_), .C(_243_), .Y(_246_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__6_), .Y(_247_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_152__bF_buf1), .C(_148__bF_buf2), .Y(_248_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__6_), .Y(_249_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_155__bF_buf2), .Y(_250_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_250_), .C(_248_), .Y(_251_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_251_), .Y(_252_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_252_), .C(_241_), .Y(AI_6_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_815__bF_buf2), .C(_1064_), .D(_125_), .Y(_253_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(ADD_7_), .C(_253_), .Y(_254_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(AXYS_1__7_), .Y(_255_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_256_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__7_), .Y(_257_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_155__bF_buf1), .Y(_258_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_258_), .C(_256_), .Y(_259_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(AXYS_3__7_), .Y(_260_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_152__bF_buf3), .C(_148__bF_buf0), .Y(_261_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__7_), .Y(_262_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_155__bF_buf0), .Y(_263_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_263_), .C(_261_), .Y(_264_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_264_), .Y(_265_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_265_), .C(_254_), .Y(AI_7_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(op_0_), .Y(_266_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_267_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_1130_), .C(_81_), .Y(_268_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_269_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf1), .B(_915_), .C(_269_), .Y(_270_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_121_), .Y(_271_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_815__bF_buf1), .B(_271_), .Y(_272_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_272_), .Y(_273_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_267_), .C(_273_), .Y(alu_op_0_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(op_1_), .Y(_274_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_267_), .C(_273_), .Y(alu_op_1_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(backwards), .Y(_275_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_276_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(op_2_), .B(_81_), .C(_276_), .Y(_277_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_815__bF_buf0), .C(_277_), .Y(alu_op_2_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(op_3_), .Y(_278_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_267_), .Y(alu_op_3_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(store), .Y(_279_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf0), .B(_1145_), .C(_271_), .Y(_280_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_280_), .Y(_281_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_1190_), .Y(_282_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_282_), .C(_281_), .Y(_1441_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .Y(_283_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(C), .B(ADD_0_), .S(php), .Y(_284_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_817_), .C(_284_), .D(_114_), .Y(_285_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_283_), .C(_285_), .Y(_286_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_287_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(PC_8_), .B(_132_), .C(PC_0_), .D(_287_), .Y(_288_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .Y(_289_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_163_), .C(_289_), .Y(_1440__0_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(php), .Y(_290_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_114_), .C(_817_), .Y(_291_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(PC_9_), .B(_132_), .C(PC_1_), .D(_287_), .Y(_292_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(php), .B(_114_), .C(_1192_), .Y(_293_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_293_), .Y(_294_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_294_), .C(_292_), .Y(_295_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(Z), .B(_291_), .C(_295_), .Y(_296_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_186_), .C(_296_), .Y(_1440__1_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_293_), .Y(_297_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_269_), .C(_956_), .D(_106_), .Y(_298_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(I), .B(_291_), .C(_298_), .Y(_299_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_297_), .Y(_300_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_199_), .C(_300_), .Y(_1440__2_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_114_), .Y(_301_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_301_), .C(D), .Y(_302_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_269_), .C(_944_), .D(_106_), .Y(_303_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_293_), .C(_303_), .Y(_304_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_302_), .Y(_305_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_212_), .C(_305_), .Y(_1440__3_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_1323_), .C(ADD_4_), .D(_301_), .Y(_306_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_829_), .C(_306_), .Y(_307_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_269_), .C(_872_), .D(_106_), .Y(_308_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_307_), .Y(_309_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_225_), .C(_309_), .Y(_1440__4_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_1323_), .C(ADD_5_), .D(_301_), .Y(_310_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_269_), .C(_817_), .Y(_311_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(PC_5_), .B(_287_), .C(_311_), .Y(_312_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_310_), .Y(_313_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_239_), .C(_313_), .Y(_1440__5_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_291_), .Y(_314_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(PC_14_), .B(_132_), .C(PC_6_), .D(_287_), .Y(_315_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_314_), .C(_315_), .Y(_316_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_293_), .C(_316_), .Y(_317_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_252_), .C(_317_), .Y(_1440__6_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(N), .Y(_318_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(PC_15_), .B(_132_), .C(PC_7_), .D(_287_), .Y(_319_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_314_), .C(_319_), .Y(_320_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_293_), .C(_320_), .Y(_321_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_265_), .C(_321_), .Y(_1440__7_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(D), .B(adc_sbc), .Y(_14_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(adc_bcd), .Y(_322_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_1205_), .Y(ALU_BCD) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_1175_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(res), .Y(_323_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_859__bF_buf0), .C(_1175_), .Y(_31_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(plp), .Y(_324_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_822__bF_buf3), .Y(_325_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_325_), .C(_169_), .Y(_326_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_325_), .C(_326_), .Y(_327_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_916_), .Y(_328_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(DIMUX_2_), .C(_328_), .Y(_329_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .Y(_330_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(sei), .Y(_331_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_331_), .C(cli), .Y(_332_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_169_), .C(_330_), .Y(_333_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_327_), .C(_329_), .Y(_6_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(shift_right), .Y(alu_shift_right) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_795__bF_buf3), .C(_916_), .Y(_334_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf2), .B(_1171_), .C(_136_), .Y(_335_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .Y(_336_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf4), .B(_1119_), .C(_1201_), .Y(_337_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(load_reg), .Y(_338_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(_338_), .Y(_339_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf3), .B(_339_), .C(_337_), .Y(_340_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_340_), .C(_1017__bF_buf5), .Y(_341_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_152__bF_buf2), .B(_341_), .C(_148__bF_buf3), .Y(_342_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_342_), .Y(_343_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf1), .B(_1171_), .C(_904_), .Y(_344_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(_43_), .C(_344_), .Y(_345_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_147_), .S(_343_), .Y(_1442__0_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(adc_bcd), .B(HC), .Y(_346_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(adj_bcd), .B(_346_), .Y(_347_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(adc_bcd), .B(adj_bcd), .C(HC), .Y(_348_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_347_), .Y(_349_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_349_), .Y(_350_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_350_), .Y(_351_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_350_), .Y(_352_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_352_), .Y(_353_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_1_), .B(_1291_), .C(_351_), .D(_353_), .Y(_354_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_176_), .S(_343_), .Y(_1442__1_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(ADD_2_), .Y(_355_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_355_), .Y(_356_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_350_), .C(_356_), .Y(_357_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_355_), .C(_1291_), .Y(_358_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_2_), .B(_1291_), .C(_357_), .D(_358_), .Y(_359_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_189_), .S(_343_), .Y(_1442__2_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .Y(_360_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_352_), .Y(_361_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_348_), .C(_361_), .Y(_362_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .Y(_363_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_363_), .Y(_364_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_364_), .Y(_365_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(DIMUX_3_), .S(_43_), .Y(_366_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_202_), .S(_343_), .Y(_1442__3_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .Y(_367_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf0), .B(_1171_), .C(_367_), .Y(_368_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_4_), .B(_43_), .C(_368_), .Y(_369_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_215_), .S(_343_), .Y(_1442__4_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(CO), .Y(_370_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(adj_bcd), .B(_370_), .C(_322_), .Y(_371_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(CO), .B(adc_bcd), .C(adj_bcd), .Y(_372_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_371_), .Y(_373_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_373_), .Y(_374_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_374_), .Y(_375_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_374_), .Y(_376_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_376_), .Y(_377_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_5_), .B(_1291_), .C(_375_), .D(_377_), .Y(_378_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_229_), .S(_343_), .Y(_1442__5_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(ADD_6_), .Y(_379_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_379_), .Y(_380_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_374_), .C(_380_), .Y(_381_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_379_), .C(_1291_), .Y(_382_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_6_), .B(_1291_), .C(_381_), .D(_382_), .Y(_383_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_242_), .S(_343_), .Y(_1442__6_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .Y(_384_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_376_), .Y(_385_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_372_), .C(_385_), .Y(_386_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .Y(_387_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_387_), .Y(_388_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_388_), .Y(_389_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(DIMUX_7_), .S(_43_), .Y(_390_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_255_), .S(_343_), .Y(_1442__7_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(NMI_1), .Y(_391_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(NMI), .B(_824_), .C(_391_), .Y(_392_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_328_), .C(_392_), .Y(_7_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(cond_code_0_), .B(_1017__bF_buf4), .Y(_393_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1361_), .C(_393_), .Y(_22__0_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(cond_code_1_), .B(_1017__bF_buf2), .Y(_394_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_1226_), .C(_394_), .Y(_22__1_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(cond_code_2_), .B(_1017__bF_buf0), .Y(_395_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf7), .B(_1090_), .C(_395_), .Y(_22__2_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_1266_), .Y(_396_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_1070__bF_buf2), .C(_1294_), .D(_396_), .Y(_30_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .Y(_397_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf2), .B(_1275_), .Y(_398_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_398_), .Y(_399_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_1070__bF_buf1), .C(_399_), .D(_397_), .Y(_29_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf6), .B(_822__bF_buf2), .C(clc), .Y(_400_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf1), .B(_1093_), .C(_1102_), .Y(_401_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_398_), .C(_1266_), .Y(_402_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_402_), .C(_400_), .Y(_17_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_822__bF_buf1), .C(sec), .Y(_403_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1361_), .Y(_404_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_404_), .Y(_405_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_402_), .C(_403_), .Y(_33_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf4), .B(_822__bF_buf0), .C(cld), .Y(_406_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_1101__bF_buf1), .Y(_407_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1226_), .Y(_408_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_1266_), .Y(_409_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_409_), .C(_406_), .Y(_18_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_822__bF_buf4), .C(sed), .Y(_410_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_404_), .Y(_411_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_409_), .C(_410_), .Y(_34_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_822__bF_buf3), .C(cli), .Y(_412_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1267_), .Y(_413_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_1266_), .Y(_414_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_414_), .C(_412_), .Y(_19_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_1070__bF_buf4), .C(_411_), .D(_414_), .Y(_35_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1275_), .Y(_415_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_404_), .Y(_416_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_822__bF_buf2), .C(clv), .Y(_417_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_396_), .C(_417_), .Y(_20_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf0), .B(_1084_), .C(_1080_), .Y(_418_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_418_), .Y(_419_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf4), .B(_1082_), .C(_419_), .Y(_420_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_1294_), .Y(_421_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_822__bF_buf1), .C(bit_ins), .Y(_422_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf0), .B(_421_), .C(_422_), .Y(_16_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1388_), .Y(_423_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_408_), .Y(_424_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .Y(_425_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1094_), .Y(_426_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .B(_426_), .C(_425_), .Y(_427_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1095_), .C(_1266_), .Y(_428_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_427_), .C(_1275_), .D(_428_), .Y(_429_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_424_), .Y(_430_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_424_), .Y(_431_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_1136_), .C(_1279_), .D(_431_), .Y(_432_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1227_), .C(_1359_), .Y(_433_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_432_), .Y(_434_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_434_), .Y(_435_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1299_), .C(_425_), .Y(_436_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_436_), .Y(_437_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_1388_), .Y(_438_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_420_), .C(_438_), .Y(_439_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_439_), .Y(_440_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_435_), .Y(_441_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_441_), .Y(_442_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_423_), .C(_442_), .Y(_443_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_444_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_420_), .Y(_445_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1358_), .C(_1070__bF_buf3), .Y(_446_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_445_), .Y(_447_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_436_), .C(_447_), .Y(_448_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_444_), .Y(_449_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_1101__bF_buf3), .C(_449_), .D(_443_), .Y(_28__0_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1183_), .Y(_450_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_1090_), .C(_446_), .Y(_451_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_451_), .Y(_452_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_1101__bF_buf2), .C(_441_), .D(_452_), .Y(_28__1_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf7), .B(_822__bF_buf0), .C(op_2_), .Y(_453_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf1), .B(_442_), .C(_453_), .Y(_28__2_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_1101__bF_buf0), .C(_436_), .D(_447_), .Y(_28__3_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1094_), .C(_419_), .Y(_454_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_454_), .Y(_455_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1359_), .C(_455_), .Y(_456_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf6), .B(_822__bF_buf4), .C(rotate), .Y(_457_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf3), .B(_456_), .C(_457_), .Y(_32_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_822__bF_buf3), .C(shift_right), .Y(_458_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf2), .B(_438_), .C(_458_), .Y(_37_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_1267_), .C(_1101__bF_buf1), .Y(_459_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_1101__bF_buf0), .C(_459_), .D(_432_), .Y(_21_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1181_), .C(_1070__bF_buf2), .Y(_460_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_1070__bF_buf1), .C(_460_), .D(_423_), .Y(_36_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf2), .B(_1123_), .C(RDY_bF_buf4), .Y(_461_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_461_), .Y(_462_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(D), .B(_1090_), .Y(_463_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1183_), .Y(_464_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_464_), .Y(_465_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_462_), .C(_463_), .D(_465_), .Y(_12_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(adc_sbc), .Y(_466_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_462_), .C(_465_), .Y(_13_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1087_), .C(_454_), .Y(_467_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_467_), .Y(_468_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf4), .B(_822__bF_buf2), .C(inc), .Y(_469_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf3), .B(_468_), .C(_469_), .Y(_24_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf3), .B(_341_), .Y(_470_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_470_), .Y(_471_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__0_), .B(_471_), .Y(_472_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_471_), .C(_472_), .Y(_1443__0_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__1_), .B(_471_), .Y(_473_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_471_), .C(_473_), .Y(_1443__1_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__2_), .B(_471_), .Y(_474_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_471_), .C(_474_), .Y(_1443__2_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__3_), .B(_471_), .Y(_475_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_471_), .C(_475_), .Y(_1443__3_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__4_), .B(_471_), .Y(_476_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_471_), .C(_476_), .Y(_1443__4_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__5_), .B(_471_), .Y(_477_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_471_), .C(_477_), .Y(_1443__5_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__6_), .B(_471_), .Y(_478_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_471_), .C(_478_), .Y(_1443__6_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(AXYS_0__7_), .B(_471_), .Y(_479_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_471_), .C(_479_), .Y(_1443__7_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_415_), .Y(_480_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_822__bF_buf1), .C(load_only), .Y(_481_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1101__bF_buf2), .B(_480_), .C(_481_), .Y(_26_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_415_), .Y(_482_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1388_), .C(_482_), .Y(_483_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1070__bF_buf0), .C(_483_), .Y(_40_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1094_), .Y(_484_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_425_), .C(_484_), .Y(_485_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_1070__bF_buf4), .C(_399_), .D(_485_), .Y(_39_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_482_), .Y(_486_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1331_), .C(_486_), .Y(_487_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(index_y), .S(_1070__bF_buf3), .Y(_488_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_488_), .C(_487_), .Y(_25_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(src_reg_0_), .Y(_489_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_426_), .C(_1086_), .Y(_490_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_482_), .Y(_491_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_491_), .Y(_492_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(_492_), .C(_490_), .Y(_493_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_825__bF_buf3), .B(_1093_), .C(_1178_), .Y(_494_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_430_), .Y(_495_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_495_), .C(_428_), .Y(_496_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_493_), .Y(_497_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_416_), .C(_497_), .Y(_498_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_498_), .Y(_499_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_1070__bF_buf1), .C(_499_), .Y(_38__0_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_1095_), .Y(_500_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_1389_), .C(_1070__bF_buf0), .Y(_501_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1077_), .Y(_502_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_502_), .C(_486_), .Y(_503_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_495_), .C(_503_), .Y(_504_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_504_), .Y(_505_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_1101__bF_buf1), .C(_505_), .D(_497_), .Y(_38__1_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(dst_reg_0_), .Y(_506_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1080_), .C(_1086_), .Y(_507_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_507_), .C(_428_), .Y(_508_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_492_), .C(_397_), .Y(_509_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_509_), .C(_1070__bF_buf4), .Y(_510_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_1070__bF_buf3), .C(_510_), .Y(_23__0_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_486_), .C(_501_), .Y(_511_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_409_), .C(_511_), .Y(_512_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_512_), .Y(_513_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_1101__bF_buf0), .C(_513_), .Y(_23__1_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_416_), .C(_433_), .Y(_514_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_416_), .Y(_515_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1085_), .Y(_516_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_415_), .C(_502_), .Y(_517_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1389_), .C(_517_), .Y(_518_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_518_), .Y(_519_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1292_), .C(_519_), .Y(_520_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_484_), .C(_1102_), .D(_1087_), .Y(_521_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_521_), .Y(_522_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_522_), .C(_1070__bF_buf2), .Y(_523_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_1070__bF_buf1), .C(_523_), .Y(_27_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1251_), .C(RDY_bF_buf3), .Y(_524_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(reset), .Y(_525_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_524_), .C(IRHOLD_0_), .Y(_526_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_525_), .C(_526_), .Y(_4__0_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_524_), .C(IRHOLD_1_), .Y(_527_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_525_), .C(_527_), .Y(_4__1_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_524_), .C(IRHOLD_2_), .Y(_528_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_525_), .C(_528_), .Y(_4__2_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_524_), .C(IRHOLD_3_), .Y(_529_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_525_), .C(_529_), .Y(_4__3_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_4_), .Y(_530_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_1019_), .S(_525_), .Y(_4__4_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_5_), .Y(_531_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_119_), .S(_525_), .Y(_4__5_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_6_), .Y(_532_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_1052_), .S(_525_), .Y(_4__6_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(IRHOLD_7_), .Y(_533_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_1064_), .S(_525_), .Y(_4__7_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_822__bF_buf0), .C(IRHOLD_valid), .Y(_534_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(reset), .B(_534_), .C(_525_), .Y(_5_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_466_), .C(plp), .Y(_535_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(AV), .C(_535_), .Y(_536_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(clv), .B(_536_), .Y(_537_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(plp), .C(_537_), .Y(_538_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(bit_ins), .Y(_539_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_1205_), .Y(_540_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_6_), .B(_540_), .Y(_541_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_540_), .C(_541_), .Y(_542_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_859__bF_buf1), .B(_1155_), .Y(_543_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_6_), .B(_1155_), .C(_543_), .D(_542_), .Y(_544_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_822__bF_buf4), .B(_538_), .C(_544_), .Y(_10_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_3_), .B(_1155_), .Y(_545_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(cld), .Y(_546_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(D), .B(sed), .C(_546_), .Y(_547_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_324_), .C(_547_), .Y(_548_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(D), .B(_548_), .S(_822__bF_buf3), .Y(_549_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_549_), .C(_545_), .Y(_3_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_470_), .Y(_550_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__0_), .B(_550_), .Y(_551_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_550_), .C(_551_), .Y(_1444__0_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__1_), .B(_550_), .Y(_552_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_550_), .C(_552_), .Y(_1444__1_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__2_), .B(_550_), .Y(_553_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_550_), .C(_553_), .Y(_1444__2_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__3_), .B(_550_), .Y(_554_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_550_), .C(_554_), .Y(_1444__3_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__4_), .B(_550_), .Y(_555_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_550_), .C(_555_), .Y(_1444__4_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__5_), .B(_550_), .Y(_556_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_550_), .C(_556_), .Y(_1444__5_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__6_), .B(_550_), .Y(_557_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_550_), .C(_557_), .Y(_1444__6_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(AXYS_2__7_), .B(_550_), .Y(_558_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_550_), .C(_558_), .Y(_1444__7_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(AN), .Y(_559_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_155__bF_buf2), .C(load_reg), .Y(_560_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_86_), .C(_559_), .Y(_561_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_560_), .Y(_562_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_562_), .C(_324_), .Y(_563_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(plp), .C(_822__bF_buf2), .Y(_564_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_563_), .C(_564_), .Y(_565_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_1205_), .C(_330_), .Y(_566_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(N), .B(_543_), .Y(_567_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_567_), .C(_1192_), .Y(_568_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_7_), .B(_566_), .C(_568_), .Y(_569_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_283_), .C(_569_), .D(_565_), .Y(_8_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(AZ), .Y(_570_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_539_), .C(_560_), .Y(_571_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(AZ), .Y(_572_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_571_), .C(_324_), .Y(_573_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(plp), .C(_822__bF_buf1), .Y(_574_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_573_), .C(_574_), .Y(_575_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_330_), .C(_1192_), .Y(_576_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(Z), .C(_576_), .Y(_577_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_283_), .C(_577_), .D(_575_), .Y(_11_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_1192_), .Y(_578_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(_466_), .Y(_579_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(plp), .B(clc), .Y(_580_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(C), .B(sec), .C(_580_), .Y(_581_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_324_), .C(_581_), .Y(_582_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(write_back), .B(_822__bF_buf0), .Y(_583_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_582_), .C(_583_), .Y(_584_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_579_), .C(_584_), .Y(_585_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_583_), .C(_330_), .Y(_586_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(DIMUX_0_), .B(_330_), .C(_586_), .D(_585_), .Y(_587_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(CO), .B(_578_), .Y(_588_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_587_), .C(_588_), .Y(_2_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_342_), .Y(_589_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_158_), .S(_589_), .Y(_1445__0_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_181_), .S(_589_), .Y(_1445__1_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_194_), .S(_589_), .Y(_1445__2_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_207_), .S(_589_), .Y(_1445__3_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_220_), .S(_589_), .Y(_1445__4_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_234_), .S(_589_), .Y(_1445__5_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_247_), .S(_589_), .Y(_1445__6_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_260_), .S(_589_), .Y(_1445__7_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(DI[7]), .Y(_590_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_275_), .C(_590_), .Y(_15_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_270_), .Y(_591_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_162_), .C(_591_), .Y(_592_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_94_), .Y(_593_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_136_), .C(_593_), .Y(_594_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_594_), .Y(_595_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf1), .B(_1071_), .C(_1211_), .Y(_596_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_91_), .Y(_597_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_911_), .Y(_598_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf4), .B(_1071_), .C(_598_), .Y(_599_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_599_), .Y(_600_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_809__bF_buf0), .B(_1138_), .C(_1109_), .Y(_601_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_795__bF_buf3), .B(_1236_), .C(_1115_), .Y(_602_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_601_), .Y(_603_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_600_), .C(_595_), .Y(_604_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf3), .B(_1145_), .C(_80_), .Y(_605_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_849__bF_buf1), .Y(_606_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_920_), .Y(_607_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_607_), .C(_1197_), .Y(_608_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_799__bF_buf2), .B(_1138_), .C(_1320_), .Y(_609_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_609_), .Y(_610_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_591_), .Y(_611_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_606_), .Y(_612_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_604_), .Y(_613_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(ABL_0_), .Y(_614_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_849__bF_buf0), .C(DIMUX_0_), .D(_609_), .Y(_615_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_605_), .Y(_616_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_0_), .C(_617_), .Y(_618_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_613_), .C(_618_), .Y(_619_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_592_), .Y(_1439__0_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_1196_), .C(_794_), .Y(_620_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_621_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_543_), .Y(_622_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_838_), .C(_1312_), .Y(_623_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_623_), .C(_598_), .Y(_624_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_624_), .Y(_625_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_870_), .Y(_626_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_164_), .Y(_627_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_627_), .Y(_628_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_628_), .Y(_629_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_625_), .C(_629_), .Y(_630_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_96_), .Y(_631_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_620_), .C(_114_), .Y(_632_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_108_), .Y(_633_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_1072_), .Y(_634_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_634_), .C(_543_), .Y(_635_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1099_), .Y(_636_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1291_), .Y(_637_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_638_), .Y(_639_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_633_), .C(_639_), .Y(_640_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_601_), .Y(_641_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_609_), .Y(_642_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_641_), .Y(_643_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1115_), .C(_1150_), .Y(_644_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_1114_), .C(_1404_), .Y(_645_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_645_), .Y(_646_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_647_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_647_), .Y(_648_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_648_), .C(_643_), .Y(_649_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_640_), .C(_649_), .Y(_650_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_650_), .Y(_651_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_592_), .C(_651__bF_buf4), .Y(_652_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_651__bF_buf3), .C(_652_), .Y(_1__0_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_185_), .C(_591_), .Y(_653_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(ABL_1_), .Y(_654_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_849__bF_buf4), .C(DIMUX_1_), .D(_609_), .Y(_655_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_616_), .C(_655_), .Y(_656_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_1_), .C(_656_), .Y(_657_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_613_), .C(_657_), .Y(_658_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_653_), .Y(_1439__1_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_653_), .C(_651__bF_buf2), .Y(_659_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_651__bF_buf1), .C(_659_), .Y(_1__1_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_198_), .C(_591_), .Y(_660_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_849__bF_buf3), .C(DIMUX_2_), .D(_609_), .Y(_661_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_616_), .C(_661_), .Y(_662_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_2_), .C(_662_), .Y(_663_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_613_), .C(_663_), .Y(_664_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_660_), .Y(_1439__2_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_660_), .C(_651__bF_buf0), .Y(_665_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_651__bF_buf4), .C(_665_), .Y(_1__2_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_211_), .C(_591_), .Y(_666_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_849__bF_buf2), .C(DIMUX_3_), .D(_609_), .Y(_667_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_616_), .C(_667_), .Y(_668_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_3_), .C(_668_), .Y(_669_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_613_), .C(_669_), .Y(_670_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_666_), .Y(_1439__3_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_666_), .C(_651__bF_buf3), .Y(_671_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_651__bF_buf2), .C(_671_), .Y(_1__3_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_224_), .C(_591_), .Y(_672_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_849__bF_buf1), .C(DIMUX_4_), .D(_609_), .Y(_673_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_616_), .C(_673_), .Y(_674_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_4_), .C(_674_), .Y(_675_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_613_), .C(_675_), .Y(_676_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_672_), .Y(_1439__4_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_672_), .C(_651__bF_buf1), .Y(_677_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_651__bF_buf0), .C(_677_), .Y(_1__4_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_238_), .C(_591_), .Y(_678_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .B(_849__bF_buf0), .C(DIMUX_5_), .D(_609_), .Y(_679_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_616_), .C(_679_), .Y(_680_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_5_), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_613_), .C(_681_), .Y(_682_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_678_), .Y(_1439__5_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_678_), .C(_651__bF_buf4), .Y(_683_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_651__bF_buf3), .C(_683_), .Y(_1__5_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_251_), .C(_591_), .Y(_684_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_849__bF_buf4), .C(DIMUX_6_), .D(_609_), .Y(_685_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_616_), .C(_685_), .Y(_686_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_6_), .C(_686_), .Y(_687_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_613_), .C(_687_), .Y(_688_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_684_), .Y(_1439__6_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_684_), .C(_651__bF_buf2), .Y(_689_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_651__bF_buf1), .C(_689_), .Y(_1__6_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_264_), .C(_591_), .Y(_690_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_849__bF_buf3), .C(DIMUX_7_), .D(_609_), .Y(_691_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_616_), .C(_691_), .Y(_692_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(ADD_7_), .C(_692_), .Y(_693_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_613_), .C(_693_), .Y(_694_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_690_), .Y(_1439__7_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_690_), .C(_651__bF_buf0), .Y(_695_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_651__bF_buf4), .C(_695_), .Y(_1__7_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_283_), .C(ABH_0_), .Y(_696_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(ADD_0_), .C(_120_), .Y(_697_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_697_), .C(_591_), .Y(_698_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_600_), .C(_595_), .Y(_699_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_699_), .Y(_700_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_613_), .C(_700_), .Y(_1439__8_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1439__8_), .B(_651__bF_buf3), .Y(_701_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_651__bF_buf2), .C(_701_), .Y(_0__0_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(_600_), .Y(_702_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_608_), .Y(_703_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf2), .B(_605_), .C(ABH_1_), .Y(_704_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_703_), .C(_704_), .Y(_705_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(DIMUX_1_), .C(_705_), .Y(_706_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_613_), .C(_706_), .Y(_1439__9_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1439__9_), .B(_651__bF_buf1), .Y(_707_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_651__bF_buf0), .C(_707_), .Y(_0__1_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf1), .B(_605_), .C(ABH_2_), .Y(_708_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_703_), .C(_708_), .Y(_709_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(DIMUX_2_), .C(_709_), .Y(_710_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_613_), .C(_710_), .Y(_1439__10_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1439__10_), .B(_651__bF_buf4), .Y(_711_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_651__bF_buf3), .C(_711_), .Y(_0__2_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf0), .B(_605_), .C(ABH_3_), .Y(_712_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_703_), .C(_712_), .Y(_713_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(DIMUX_3_), .C(_713_), .Y(_714_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_613_), .C(_714_), .Y(_1439__11_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1439__11_), .B(_651__bF_buf2), .Y(_715_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_651__bF_buf1), .C(_715_), .Y(_0__3_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_703_), .C(_1019_), .D(_600_), .Y(_716_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(ABH_4_), .B(_606_), .C(_716_), .Y(_717_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_613_), .C(_717_), .Y(_1439__12_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1439__12_), .B(_651__bF_buf0), .Y(_718_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_651__bF_buf4), .C(_718_), .Y(_0__4_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf4), .B(_605_), .C(ABH_5_), .Y(_719_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_703_), .C(_719_), .Y(_720_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(DIMUX_5_), .C(_720_), .Y(_721_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_613_), .C(_721_), .Y(_1439__13_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1439__13_), .B(_651__bF_buf3), .Y(_722_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_651__bF_buf2), .C(_722_), .Y(_0__5_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(PC_14_), .Y(_723_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_849__bF_buf3), .B(_605_), .C(ABH_6_), .Y(_724_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_703_), .C(_724_), .Y(_725_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(DIMUX_6_), .C(_725_), .Y(_726_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_613_), .C(_726_), .Y(_1439__14_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1439__14_), .B(_651__bF_buf1), .Y(_727_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_651__bF_buf0), .C(_727_), .Y(_0__6_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_703_), .C(_1064_), .D(_600_), .Y(_728_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(ABH_7_), .B(_606_), .C(_728_), .Y(_729_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_613_), .C(_729_), .Y(_1439__15_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1439__15_), .B(_651__bF_buf4), .Y(_730_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_651__bF_buf3), .C(_730_), .Y(_0__7_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_820_), .C(_910_), .Y(_731_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_927_), .Y(_732_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_731_), .Y(_733_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_734_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_808_), .C(_909_), .Y(_735_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_734_), .C(_732_), .Y(_736_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_736_), .Y(_737_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_905_), .C(_733_), .D(_737_), .Y(_9__0_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_928_), .Y(_738_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_1031_), .Y(_739_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_933_), .C(_738_), .D(_739_), .Y(_9__1_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_740_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_820_), .C(_962_), .Y(_741_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_740_), .Y(_742_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_741_), .C(_928_), .Y(_743_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_743_), .Y(_744_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf4), .B(_956_), .C(_744_), .D(_742_), .Y(_9__2_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1032_), .Y(_745_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_745_), .Y(_746_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_743_), .C(RDY_bF_buf3), .Y(_747_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf2), .B(_944_), .C(_746_), .D(_747_), .Y(_9__3_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_820_), .C(_878_), .Y(_748_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_743_), .Y(_749_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_748_), .C(_1017__bF_buf0), .Y(_750_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_749_), .C(_750_), .Y(_751_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_872_), .C(_751_), .Y(_9__4_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_820_), .C(_867_), .Y(_752_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_748_), .C(_752_), .Y(_753_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_754_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_754_), .C(_743_), .Y(_755_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_1017__bF_buf7), .Y(_756_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf0), .B(_860_), .C(_753_), .D(_756_), .Y(_9__5_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_820_), .C(_899_), .Y(_757_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_757_), .C(_1017__bF_buf6), .Y(_758_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_755_), .C(_758_), .Y(_759_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_893_), .C(_759_), .Y(_9__6_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_820_), .C(_889_), .Y(_760_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_757_), .C(_760_), .Y(_761_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_757_), .C(_755_), .Y(_762_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf7), .B(_762_), .Y(_763_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_883_), .C(_761_), .D(_763_), .Y(_9__7_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_820_), .C(_1012_), .Y(_764_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_964_), .C(_764_), .Y(_765_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_1030_), .C(_740_), .Y(_766_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_764_), .Y(_767_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .B(_765_), .C(_767_), .Y(_768_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf5), .B(_1008_), .Y(_769_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_769_), .Y(_9__8_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_820_), .C(_1000_), .Y(_770_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_964_), .Y(_771_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_764_), .C(_770_), .Y(_772_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .Y(_773_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_766_), .C(RDY_bF_buf4), .Y(_774_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf3), .B(_996_), .C(_772_), .D(_774_), .Y(_9__9_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_820_), .C(_987_), .Y(_775_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_766_), .Y(_776_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_776_), .Y(_777_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_775_), .Y(_778_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_771_), .Y(_779_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_779_), .C(RDY_bF_buf2), .Y(_780_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf1), .B(_983_), .C(_780_), .D(_777_), .Y(_9__10_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_820_), .C(_976_), .Y(_781_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_776_), .B(_775_), .C(_781_), .Y(_782_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_766_), .C(RDY_bF_buf0), .Y(_783_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf8), .B(_972_), .C(_783_), .D(_782_), .Y(_9__11_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1015_), .Y(_784_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .Y(_785_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1043_), .C(RDY_bF_buf7), .Y(_786_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf6), .B(_1016_), .C(_784_), .D(_786_), .Y(_9__12_) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1439__0_), .Y(AB[0]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_1439__1_), .Y(AB[1]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_1439__2_), .Y(AB[2]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_1439__3_), .Y(AB[3]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1439__4_), .Y(AB[4]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_1439__5_), .Y(AB[5]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1439__6_), .Y(AB[6]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1439__7_), .Y(AB[7]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1439__8_), .Y(AB[8]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1439__9_), .Y(AB[9]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1439__10_), .Y(AB[10]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1439__11_), .Y(AB[11]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1439__12_), .Y(AB[12]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1439__13_), .Y(AB[13]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_1439__14_), .Y(AB[14]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_1439__15_), .Y(AB[15]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1440__0_), .Y(DO[0]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_1440__1_), .Y(DO[1]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_1440__2_), .Y(DO[2]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_1440__3_), .Y(DO[3]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_1440__4_), .Y(DO[4]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_1440__5_), .Y(DO[5]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_1440__6_), .Y(DO[6]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_1440__7_), .Y(DO[7]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .Y(WE) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1443__0_), .Q(AXYS_0__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1443__1_), .Q(AXYS_0__1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1443__2_), .Q(AXYS_0__2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1443__3_), .Q(AXYS_0__3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1443__4_), .Q(AXYS_0__4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1443__5_), .Q(AXYS_0__5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1443__6_), .Q(AXYS_0__6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1443__7_), .Q(AXYS_0__7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1442__0_), .Q(AXYS_1__0_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1442__1_), .Q(AXYS_1__1_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1442__2_), .Q(AXYS_1__2_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1442__3_), .Q(AXYS_1__3_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1442__4_), .Q(AXYS_1__4_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1442__5_), .Q(AXYS_1__5_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1442__6_), .Q(AXYS_1__6_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1442__7_), .Q(AXYS_1__7_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1445__0_), .Q(AXYS_3__0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1445__1_), .Q(AXYS_3__1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1445__2_), .Q(AXYS_3__2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1445__3_), .Q(AXYS_3__3_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1445__4_), .Q(AXYS_3__4_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1445__5_), .Q(AXYS_3__5_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1445__6_), .Q(AXYS_3__6_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1445__7_), .Q(AXYS_3__7_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1444__0_), .Q(AXYS_2__0_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1444__1_), .Q(AXYS_2__1_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1444__2_), .Q(AXYS_2__2_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1444__3_), .Q(AXYS_2__3_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1444__4_), .Q(AXYS_2__4_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1444__5_), .Q(AXYS_2__5_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1444__6_), .Q(AXYS_2__6_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1444__7_), .Q(AXYS_2__7_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_7_), .Q(NMI_edge) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(NMI), .Q(NMI_1) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_22__0_), .Q(cond_code_0_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_22__1_), .Q(cond_code_1_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_22__2_), .Q(cond_code_2_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_30_), .Q(plp) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_29_), .Q(php) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17_), .Q(clc) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_33_), .Q(sec) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_18_), .Q(cld) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_34_), .Q(sed) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_19_), .Q(cli) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_35_), .Q(sei) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20_), .Q(clv) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_16_), .Q(bit_ins) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_28__0_), .Q(op_0_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_28__1_), .Q(op_1_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_28__2_), .Q(op_2_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_28__3_), .Q(op_3_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_32_), .Q(rotate) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_37_), .Q(shift_right) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21_), .Q(compare) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_36_), .Q(shift) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_12_), .Q(adc_bcd) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_13_), .Q(adc_sbc) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_24_), .Q(inc) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_26_), .Q(load_only) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_40_), .Q(write_back) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_39_), .Q(store) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_25_), .Q(index_y) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_38__0_), .Q(src_reg_0_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_38__1_), .Q(src_reg_1_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_23__0_), .Q(dst_reg_0_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_23__1_), .Q(dst_reg_1_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_27_), .Q(load_reg) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_31_), .Q(res) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(DIMUX_0_), .Q(DIHOLD_0_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(DIMUX_1_), .Q(DIHOLD_1_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(DIMUX_2_), .Q(DIHOLD_2_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(DIMUX_3_), .Q(DIHOLD_3_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(DIMUX_4_), .Q(DIHOLD_4_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(DIMUX_5_), .Q(DIHOLD_5_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(DIMUX_6_), .Q(DIHOLD_6_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(DIMUX_7_), .Q(DIHOLD_7_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_4__0_), .Q(IRHOLD_0_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_4__1_), .Q(IRHOLD_1_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_4__2_), .Q(IRHOLD_2_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_4__3_), .Q(IRHOLD_3_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4__4_), .Q(IRHOLD_4_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4__5_), .Q(IRHOLD_5_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4__6_), .Q(IRHOLD_6_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_4__7_), .Q(IRHOLD_7_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_5_), .Q(IRHOLD_valid) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_10_), .Q(V) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3_), .Q(D) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_6_), .Q(I) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_8_), .Q(N) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_11_), .Q(Z) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2_), .Q(C) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_15_), .Q(backwards) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_14_), .Q(adj_bcd) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1__0_), .Q(ABL_0_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1__1_), .Q(ABL_1_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1__2_), .Q(ABL_2_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1__3_), .Q(ABL_3_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1__4_), .Q(ABL_4_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1__5_), .Q(ABL_5_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1__6_), .Q(ABL_6_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1__7_), .Q(ABL_7_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__0_), .Q(ABH_0_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__1_), .Q(ABH_1_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__2_), .Q(ABH_2_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__3_), .Q(ABH_3_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__4_), .Q(ABH_4_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__5_), .Q(ABH_5_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__6_), .Q(ABH_6_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_0__7_), .Q(ABH_7_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_9__0_), .Q(PC_0_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_9__1_), .Q(PC_1_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_9__2_), .Q(PC_2_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_9__3_), .Q(PC_3_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_9__4_), .Q(PC_4_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__5_), .Q(PC_5_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_9__6_), .Q(PC_6_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_9__7_), .Q(PC_7_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_9__8_), .Q(PC_8_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_9__9_), .Q(PC_9_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_9__10_), .Q(PC_10_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__11_), .Q(PC_11_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_9__12_), .Q(PC_12_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_9__13_), .Q(PC_13_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_9__14_), .Q(PC_14_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_9__15_), .Q(PC_15_) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1438__0_), .Q(state_0_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1438__1_), .Q(state_1_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1438__2_), .Q(state_2_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1438__3_), .Q(state_3_), .R(vdd), .S(_1175_) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1438__4_), .Q(state_4_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1438__5_), .Q(state_5_), .R(_1175_), .S(vdd) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(ADD_0_), .Y(_1626_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(ADD_7_), .Y(_1627_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(ADD_5_), .Y(_1628_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(ADD_1_), .Y(_1629_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_1628_), .C(_1629_), .Y(_1630_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .B(_1630_), .Y(AZ) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(RDY_bF_buf5), .Y(_1631_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(CO), .B(_1631__bF_buf3), .Y(_1632_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(alu_op_3_), .Y(_1633_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(_1633_), .Y(_1634_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .Y(_1635_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(alu_op_1_), .B(_1635_), .Y(_1636_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(BI_5_), .Y(_1637_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1637_), .Y(_1638_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(alu_op_1_), .Y(_1639_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(AI_5_), .Y(_1640_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1640_), .C(BI_5_), .Y(_1641_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1638_), .C(_1641_), .Y(_1642_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(_1638_), .Y(_1643_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1640_), .C(alu_shift_right), .Y(_1644_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(AI_6_), .C(_1642_), .D(_1644_), .Y(_1645_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .Y(_1646_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .Y(_1647_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(alu_op_3_), .B(_1647_), .Y(_1648_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_5_), .Y(_1649_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(BI_5_), .B(_1648_), .C(_1649_), .Y(_1650_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .Y(_1651_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1651_), .C(_1646_), .Y(_1652_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .Y(_1653_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .Y(_1654_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1639_), .Y(_1655_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(BI_4_), .Y(_1656_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(AI_4_), .B(_1656_), .Y(_1657_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(BI_4_), .C(_1655_), .D(_1657_), .Y(_1658_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(AI_4_), .B(_1656_), .C(_1654_), .Y(_1659_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1640_), .C(_1659_), .D(_1658_), .Y(_1660_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_4_), .Y(_1661_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(BI_4_), .B(_1648_), .C(_1661_), .Y(_1662_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_1662_), .Y(_1663_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1663_), .C(_1660_), .Y(_1664_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(AI_3_), .Y(_1665_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(BI_2_), .Y(_1666_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1666_), .Y(_1667_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(AI_2_), .Y(_1668_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1668_), .C(BI_2_), .Y(_1669_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1667_), .C(_1669_), .Y(_1670_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1666_), .C(_1668_), .Y(_1671_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1671_), .C(_1670_), .Y(_1452_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1665_), .C(_1452_), .Y(_1453_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_2_), .Y(_1454_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(BI_2_), .B(_1648_), .C(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(_1633_), .C(_1455_), .Y(_1456_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(AI_1_), .B(BI_1_), .C(_1635_), .Y(_1457_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(BI_1_), .C(_1655_), .D(_1457_), .Y(_1458_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(AI_1_), .Y(_1459_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(BI_1_), .Y(_1460_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1460_), .C(_1459_), .Y(_1461_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1461_), .Y(_1462_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1668_), .C(_1462_), .D(_1458_), .Y(_1463_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_1_), .Y(_1464_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(BI_1_), .B(_1648_), .C(_1464_), .Y(_1465_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .Y(_1466_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1466_), .C(_1463_), .Y(_1467_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(AI_1_), .Y(_1468_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(BI_0_), .B(_1635_), .Y(_1469_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(alu_op_1_), .B(AI_0_), .Y(_1470_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(BI_0_), .B(_1470_), .C(_1655_), .D(_1469_), .Y(_1471_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(AI_0_), .Y(_1472_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(BI_0_), .Y(_1473_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1473_), .C(_1472_), .Y(_1474_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1474_), .Y(_1475_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1475_), .C(_1468_), .Y(_1476_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_0_), .Y(_1477_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(BI_0_), .B(_1648_), .C(_1477_), .Y(_1478_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(_1633_), .C(_1478_), .Y(_1479_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_1633_), .C(CI), .Y(_1480_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(_1480_), .Y(_1481_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(alu_op_1_), .B(_1473_), .S(alu_op_0_), .Y(_1482_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(BI_0_), .B(_1470_), .Y(_1483_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1482_), .Y(_1484_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1472_), .C(alu_shift_right), .Y(_1485_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_1484_), .Y(_1486_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1478_), .C(_1486_), .Y(_1487_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_1479_), .C(_1481_), .D(_1487_), .Y(_1488_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1463_), .Y(_1489_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .B(_1488_), .C(_1467_), .Y(_1490_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(_1455_), .S(_1453_), .Y(_1491_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1456_), .C(_1491_), .D(_1490_), .Y(_1492_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(AI_4_), .Y(_1493_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(BI_3_), .Y(_1494_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1494_), .Y(_1495_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(AI_3_), .B(_1495_), .Y(_1496_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(BI_3_), .C(_1655_), .D(_1496_), .Y(_1497_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(AI_3_), .B(_1495_), .C(_1654_), .Y(_1498_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1498_), .B(_1497_), .C(_1493_), .Y(_1499_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(alu_op_3_), .B(_1647_), .C(_1494_), .Y(_1500_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_3_), .Y(_1501_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1501_), .Y(_1502_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1502_), .C(_1499_), .Y(_1503_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .B(_1502_), .C(_1503_), .Y(_1504_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1504_), .Y(_1505_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(ALU_BCD), .Y(_1506_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .Y(_1507_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1507_), .C(_1476_), .Y(_1508_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .Y(_1509_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1476_), .Y(_1510_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .B(_1510_), .C(_1508_), .Y(_1511_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(_1633_), .C(_1465_), .Y(_1512_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1512_), .C(_1489_), .Y(_1513_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1511_), .Y(_1514_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1466_), .C(_1467_), .Y(_1515_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1515_), .Y(_1516_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1514_), .Y(_1517_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1490_), .Y(_1518_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_1455_), .Y(_1519_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1519_), .C(_1453_), .Y(_1520_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1519_), .C(_1520_), .Y(_1521_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_1521_), .C(_1514_), .Y(_1522_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .B(_1522_), .Y(_1523_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1517_), .C(_1506_), .Y(_1524_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_1492_), .C(_1503_), .Y(_1525_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1505_), .C(_1525_), .Y(_1526_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1663_), .C(_1664_), .Y(_1527_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1526_), .C(_1664_), .Y(_1528_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1651_), .C(_1652_), .Y(_1529_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .Y(_1530_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1530_), .C(_1653_), .Y(_1531_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(BI_7_), .Y(_1532_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1532_), .Y(_1533_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(AI_7_), .Y(_1534_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1534_), .C(BI_7_), .Y(_1535_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1533_), .C(_1535_), .Y(_1536_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .Y(_1537_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1534_), .C(alu_shift_right), .Y(_1538_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(CI), .B(alu_shift_right), .C(_1536_), .D(_1538_), .Y(_1539_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .Y(_1540_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_7_), .Y(_1541_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(BI_7_), .B(_1648_), .C(_1541_), .Y(_1542_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .Y(_1543_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(_1634_), .C(_1540_), .Y(_1544_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .Y(_1545_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(BI_6_), .Y(_1546_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(alu_op_0_), .B(_1546_), .Y(_1547_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(AI_6_), .Y(_1548_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1548_), .C(BI_6_), .Y(_1549_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1547_), .C(_1549_), .Y(_1550_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .Y(_1551_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1548_), .C(alu_shift_right), .Y(_1552_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(AI_7_), .B(alu_shift_right), .C(_1550_), .D(_1552_), .Y(_1553_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .Y(_1554_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(alu_op_3_), .C(BI_6_), .Y(_1555_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(BI_6_), .B(_1648_), .C(_1555_), .Y(_1556_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_1556_), .Y(_1557_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1557_), .C(_1554_), .Y(_1558_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .Y(_1559_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1540_), .B(_1543_), .C(_1544_), .Y(_1560_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .Y(_1561_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1559_), .C(_1545_), .Y(_1562_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1557_), .C(_1558_), .Y(_1563_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .Y(_1564_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1561_), .Y(_1565_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1531_), .C(_1562_), .Y(_1566_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(AI_0_), .C(_1566_), .Y(_1567_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(alu_shift_right), .B(AI_0_), .Y(_1568_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1565_), .Y(_1569_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_1562_), .C(_1569_), .Y(_1570_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .Y(_1571_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1524_), .Y(_1572_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1573_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .Y(_1574_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .Y(_1575_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1575_), .B(_1574_), .C(_1662_), .Y(_1576_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .B(_1574_), .Y(_1577_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1576_), .Y(_1578_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1578_), .C(_1573_), .D(_1572_), .Y(_1579_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1579_), .C(_1530_), .Y(_1580_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1575_), .B(_1553_), .C(_1556_), .Y(_1581_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_1553_), .Y(_1582_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1581_), .Y(_1583_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1583_), .C(_1652_), .D(_1580_), .Y(_1584_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1584_), .C(_1560_), .Y(_1585_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(alu_op_2_), .B(_1633_), .C(_1662_), .Y(_1586_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1504_), .Y(_1587_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_1491_), .C(_1514_), .Y(_1588_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1490_), .Y(_1589_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(_1517_), .C(_1588_), .Y(_1590_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(ALU_BCD), .B(_1590_), .Y(_1591_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1591_), .B(_1587_), .C(_1573_), .Y(_1592_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .Y(_1593_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1586_), .C(_1593_), .D(_1592_), .Y(_1594_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1594_), .C(_1652_), .Y(_1595_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1595_), .Y(_1596_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1561_), .C(_1596_), .Y(_1597_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1585_), .Y(_1598_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1594_), .Y(_1599_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_1580_), .Y(_1600_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1563_), .C(_1580_), .Y(_1601_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1596_), .Y(_1602_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1600_), .C(_1506_), .Y(_1603_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1570_), .C(_1598_), .D(_1603_), .Y(_1604_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_1604_), .C(_1632_), .Y(_1448_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .Y(_1605_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(AN), .B(_1631__bF_buf1), .Y(_1606_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1605_), .C(_1606_), .Y(_1450_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(HC), .B(_1631__bF_buf3), .Y(_1607_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_1526_), .C(_1607_), .Y(_1449_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(ADD_0_), .B(_1631__bF_buf1), .Y(_1608_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1487_), .C(_1481_), .Y(_1609_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_1507_), .C(_1508_), .Y(_1610_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .B(_1610_), .C(RDY_bF_buf4), .Y(_1611_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1611_), .C(_1608_), .Y(_1451__0_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(ADD_1_), .B(_1631__bF_buf0), .Y(_1612_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_1517_), .C(_1612_), .Y(_1451__1_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(ADD_2_), .B(_1631__bF_buf2), .Y(_1613_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_1523_), .C(_1613_), .Y(_1451__2_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(ADD_3_), .B(_1631__bF_buf0), .Y(_1614_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_1587_), .C(_1614_), .Y(_1451__3_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(ADD_4_), .B(_1631__bF_buf2), .Y(_1615_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1592_), .Y(_1616_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1526_), .C(RDY_bF_buf3), .Y(_1617_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1617_), .C(_1615_), .Y(_1451__4_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(ADD_5_), .B(_1631__bF_buf1), .Y(_1618_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1600_), .C(_1618_), .Y(_1451__5_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(ADD_6_), .B(_1631__bF_buf3), .Y(_1619_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_1602_), .C(_1619_), .Y(_1451__6_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(ADD_7_), .B(_1631__bF_buf1), .Y(_1620_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1605_), .C(_1620_), .Y(_1451__7_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1540_), .B(_1634_), .C(_1543_), .Y(_1621_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI7), .B(_1631__bF_buf3), .Y(_1622_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_1621_), .C(_1622_), .Y(_1447_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(ALU_AI7), .B(_1631__bF_buf1), .Y(_1623_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_1534_), .B(_1631__bF_buf0), .C(_1623_), .Y(_1446_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ALU_BI7), .B(ALU_AI7), .Y(_1624_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(CO), .B(AN), .Y(_1625_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1624_), .B(_1625_), .Y(AV) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1448_), .Q(CO) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1450_), .Q(AN) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1449_), .Q(HC) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1451__0_), .Q(ADD_0_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1451__1_), .Q(ADD_1_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1451__2_), .Q(ADD_2_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1451__3_), .Q(ADD_3_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1451__4_), .Q(ADD_4_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1451__5_), .Q(ADD_5_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1451__6_), .Q(ADD_6_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1451__7_), .Q(ADD_7_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1447_), .Q(ALU_BI7) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1446_), .Q(ALU_AI7) );
endmodule
