module fp_divider ( gnd, vdd, input_a, input_b, input_a_stb, input_b_stb, output_z_ack, clk, rst, output_z, output_z_stb, input_a_ack, input_b_ack);

input gnd, vdd;
input input_a_stb;
input input_b_stb;
input output_z_ack;
input clk;
input rst;
output output_z_stb;
output input_a_ack;
output input_b_ack;
input [31:0] input_a;
input [31:0] input_b;
output [31:0] output_z;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(state_12_), .Y(state_12_bF_buf4) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(state_12_), .Y(state_12_bF_buf3) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(state_12_), .Y(state_12_bF_buf2) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(state_12_), .Y(state_12_bF_buf1) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(state_12_), .Y(state_12_bF_buf0) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_124__bF_buf3) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_124__bF_buf2) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_124__bF_buf1) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_124__bF_buf0) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_194__bF_buf3) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_194__bF_buf2) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_194__bF_buf1) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_194__bF_buf0) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf6) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf5) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf4) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf3) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf2) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf1) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf0) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf6) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf5) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf4) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf3) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf2) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf1) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(state_4_bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf56) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf55) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf54) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf52) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf51) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf50) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf49) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf48) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf46) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf45) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf44) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf43) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf42) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf41) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf40) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf39) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf38) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf37) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf36) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf35) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf34) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf33) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf32) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf31) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf30) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf29) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf26) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf25) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf24) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf23) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf22) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf21) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf20) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf19) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf18) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf17) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf15) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf14) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf13) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf12) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf11) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf10) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf9) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf8) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf7) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf6) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf5) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf4) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf3) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf2) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf1) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf0) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf6) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf5) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf4) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf3) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf2) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf1) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(state_1_bF_buf0) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf5) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf4) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf3) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf2) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf1) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_567__bF_buf0) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_36__bF_buf4) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_36__bF_buf3) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_36__bF_buf2) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_36__bF_buf1) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_36__bF_buf0) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf6) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf5) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf4) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf3) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf2) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf1) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_182__bF_buf0) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_561_), .Y(_561__bF_buf4) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_561_), .Y(_561__bF_buf3) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_561_), .Y(_561__bF_buf2) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_561_), .Y(_561__bF_buf1) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_561_), .Y(_561__bF_buf0) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .Y(_1973__bF_buf3) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .Y(_1973__bF_buf2) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .Y(_1973__bF_buf1) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .Y(_1973__bF_buf0) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf7) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf6) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf5) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf4) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf3) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf2) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf1) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(state_14_), .Y(state_14_bF_buf0) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(state_11_), .Y(state_11_bF_buf4) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(state_11_), .Y(state_11_bF_buf3) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(state_11_), .Y(state_11_bF_buf2) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(state_11_), .Y(state_11_bF_buf1) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(state_11_), .Y(state_11_bF_buf0) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf6) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf5) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf4) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf3) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf2) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf1) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_199__bF_buf0) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf7) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf6) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf5) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf4) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf3) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf2) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf1) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(state_6_bF_buf0) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(state_3_bF_buf4) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(state_3_bF_buf3) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(state_3_bF_buf2) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(state_3_bF_buf1) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(state_3_bF_buf0) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_38__bF_buf4) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_38__bF_buf3) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_38__bF_buf2) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_38__bF_buf1) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_38__bF_buf0) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf3) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf2) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf1) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf0) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf7) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf6) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf5) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf4) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf3) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf2) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf1) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_202__bF_buf0) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf6) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf5) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf4) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf3) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf2) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf1) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_563_), .Y(_563__bF_buf0) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_237__bF_buf3) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_237__bF_buf2) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_237__bF_buf1) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_237__bF_buf0) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_234__bF_buf4) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_234__bF_buf3) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_234__bF_buf2) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_234__bF_buf1) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_234__bF_buf0) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_228__bF_buf3) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_228__bF_buf2) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_228__bF_buf1) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_228__bF_buf0) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf5) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf4) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf3) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf2) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf1) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1258__bF_buf0) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf7) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf6) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf5) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf4) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf3) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf2) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf1) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(_871_), .Y(_871__bF_buf0) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf7) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf6) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf5) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf4) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf3) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf2) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf1) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_245__bF_buf0) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_239__bF_buf3) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_239__bF_buf2) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_239__bF_buf1) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_239__bF_buf0) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf6) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf5) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf4) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf3) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf2) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf1) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_562__bF_buf0) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .Y(_1974__bF_buf3) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .Y(_1974__bF_buf2) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .Y(_1974__bF_buf1) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .Y(_1974__bF_buf0) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf3) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf2) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf1) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf0) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(a_m_3_), .Y(_1968_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_4_bF_buf6), .Y(_1969_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(a_m_23_), .Y(_1970_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_1971_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_1971_), .Y(_1972_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1972_), .Y(_1973_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(a_m_23_), .B(_1971_), .Y(_1974_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(a_3_), .B(state_4_bF_buf4), .C(a_m_2_), .D(_1974__bF_buf3), .Y(_1975_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1968_), .B(_1973__bF_buf3), .C(_1975_), .Y(_2__3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(a_m_4_), .Y(_1976_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_4_), .C(a_m_3_), .D(_1974__bF_buf3), .Y(_1977_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_1973__bF_buf2), .C(_1977_), .Y(_2__4_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(a_m_5_), .Y(_1978_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_5_), .C(a_m_4_), .D(_1974__bF_buf0), .Y(_1979_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1973__bF_buf2), .C(_1979_), .Y(_2__5_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(a_m_6_), .Y(_1980_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_6_), .C(a_m_5_), .D(_1974__bF_buf0), .Y(_1981_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_1973__bF_buf2), .C(_1981_), .Y(_2__6_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(a_m_7_), .Y(_1982_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_7_), .C(a_m_6_), .D(_1974__bF_buf2), .Y(_1983_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1973__bF_buf1), .C(_1983_), .Y(_2__7_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(a_m_8_), .Y(_1984_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_8_), .C(a_m_7_), .D(_1974__bF_buf2), .Y(_1985_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1984_), .B(_1973__bF_buf1), .C(_1985_), .Y(_2__8_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(a_m_9_), .Y(_1986_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_9_), .C(a_m_8_), .D(_1974__bF_buf2), .Y(_1987_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1973__bF_buf1), .C(_1987_), .Y(_2__9_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(a_m_10_), .Y(_1988_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_10_), .C(a_m_9_), .D(_1974__bF_buf3), .Y(_1989_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1988_), .B(_1973__bF_buf3), .C(_1989_), .Y(_2__10_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(a_m_11_), .Y(_1990_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_11_), .C(a_m_10_), .D(_1974__bF_buf1), .Y(_1991_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1973__bF_buf3), .C(_1991_), .Y(_2__11_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(a_m_12_), .Y(_1992_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_12_), .C(a_m_11_), .D(_1974__bF_buf1), .Y(_1993_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_1973__bF_buf0), .C(_1993_), .Y(_2__12_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(a_m_13_), .Y(_1994_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_13_), .C(a_m_12_), .D(_1974__bF_buf1), .Y(_1995_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(_1973__bF_buf0), .C(_1995_), .Y(_2__13_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(a_m_14_), .Y(_1996_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_14_), .C(a_m_13_), .D(_1974__bF_buf1), .Y(_1997_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_1973__bF_buf0), .C(_1997_), .Y(_2__14_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(a_m_15_), .Y(_1998_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_15_), .C(a_m_14_), .D(_1974__bF_buf1), .Y(_1999_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_1973__bF_buf0), .C(_1999_), .Y(_2__15_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(a_m_16_), .Y(_2000_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_16_), .C(a_m_15_), .D(_1974__bF_buf1), .Y(_2001_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .B(_1973__bF_buf3), .C(_2001_), .Y(_2__16_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(a_m_17_), .Y(_2002_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_17_), .C(a_m_16_), .D(_1974__bF_buf2), .Y(_2003_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_1973__bF_buf3), .C(_2003_), .Y(_2__17_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(a_m_18_), .Y(_24_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_18_), .C(a_m_17_), .D(_1974__bF_buf3), .Y(_25_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_1973__bF_buf3), .C(_25_), .Y(_2__18_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(a_m_19_), .Y(_26_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf1), .B(a_19_), .C(a_m_18_), .D(_1974__bF_buf3), .Y(_27_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_1973__bF_buf1), .C(_27_), .Y(_2__19_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(a_m_20_), .Y(_28_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_20_), .C(a_m_19_), .D(_1974__bF_buf2), .Y(_29_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_1973__bF_buf1), .C(_29_), .Y(_2__20_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(a_m_21_), .Y(_30_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_21_), .C(a_m_20_), .D(_1974__bF_buf2), .Y(_31_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_1973__bF_buf2), .C(_31_), .Y(_2__21_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(a_m_22_), .Y(_32_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_22_), .C(a_m_21_), .D(_1974__bF_buf0), .Y(_33_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_1973__bF_buf2), .C(_33_), .Y(_2__22_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(z_e_9_), .Y(_34_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(z_e_8_), .B(z_e_7_), .C(_34_), .Y(_35_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_0_), .Y(_37_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf1), .B(state_11_bF_buf0), .Y(_38_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(b_e_5_), .B(b_e_4_), .Y(_39_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(b_e_6_), .Y(_41_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(b_e_7_), .B(_41_), .Y(_42_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_40_), .Y(_43_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(b_e_3_), .B(b_e_2_), .Y(_45_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(b_e_9_), .Y(_46_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(_46_), .Y(_47_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(b_e_0_), .B(b_e_8_), .Y(_48_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_47_), .C(_48_), .Y(_49_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_44_), .Y(_50_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(_51_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(b_m_21_), .Y(_52_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(b_m_20_), .Y(_53_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(b_m_23_), .B(b_m_22_), .Y(_54_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .C(_54_), .Y(_55_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(b_m_17_), .Y(_56_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(b_m_16_), .Y(_57_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(b_m_19_), .B(b_m_18_), .Y(_58_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_57_), .C(_58_), .Y(_59_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_59_), .Y(_60_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(b_m_1_), .Y(_61_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(b_m_0_), .Y(_62_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(b_m_3_), .B(b_m_2_), .Y(_63_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_62_), .C(_63_), .Y(_64_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(b_m_7_), .Y(_65_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(b_m_6_), .Y(_66_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(b_m_5_), .B(b_m_4_), .Y(_67_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(_67_), .Y(_68_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_68_), .Y(_69_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(b_m_15_), .Y(_70_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(b_m_14_), .Y(_71_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(b_m_13_), .B(b_m_12_), .Y(_72_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .C(_72_), .Y(_73_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(b_m_9_), .Y(_74_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(b_m_8_), .Y(_75_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(b_m_11_), .B(b_m_10_), .Y(_76_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_76_), .Y(_77_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_77_), .Y(_78_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_69_), .C(_78_), .Y(_79_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_51_), .C(state_12_bF_buf2), .Y(_80_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(a_e_5_), .B(a_e_4_), .Y(_81_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_82_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(a_e_6_), .Y(_83_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(a_e_7_), .B(_83_), .Y(_84_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_82_), .Y(_85_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .Y(_87_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(a_e_3_), .B(a_e_2_), .Y(_88_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(a_e_0_), .C(_88_), .Y(_89_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_86_), .Y(_90_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(a_e_9_), .B(a_e_8_), .C(_90_), .Y(_91_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(a_m_4_), .B(a_m_5_), .Y(_92_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_1982_), .C(_92_), .Y(_93_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(a_m_2_), .Y(_94_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_1968_), .Y(_95_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_32_), .Y(_96_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_96_), .Y(_97_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_97_), .Y(_98_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(a_m_12_), .B(a_m_13_), .Y(_99_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_1998_), .C(_99_), .Y(_100_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(a_m_8_), .B(a_m_9_), .Y(_101_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1988_), .B(_1990_), .C(_101_), .Y(_102_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .Y(_103_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(a_m_16_), .B(a_m_17_), .Y(_104_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_26_), .C(_104_), .Y(_105_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(a_m_1_), .B(a_m_0_), .Y(_106_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_30_), .C(_106_), .Y(_107_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_105_), .Y(_108_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_108_), .C(_98_), .Y(_109_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(a_e_9_), .Y(_110_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(a_e_8_), .Y(_111_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(a_e_0_), .Y(_112_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_112_), .Y(_113_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_113_), .Y(_114_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .Y(_115_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(b_e_0_), .Y(_116_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .C(_45_), .Y(_117_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(b_e_9_), .B(b_e_8_), .Y(_119_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_118_), .C(_43_), .Y(_120_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_86_), .C(_120_), .Y(_121_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_91_), .C(_122_), .Y(_123_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_123_), .Y(_124_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_0_), .Y(_125_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_37_), .C(_125_), .Y(_20__0_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_1_), .Y(_126_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_1_), .Y(_127_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_126_), .C(_127_), .Y(_20__1_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_2_), .Y(_128_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf2), .B(_124__bF_buf1), .C(z_2_), .Y(_129_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_128_), .C(_129_), .Y(_20__2_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_3_), .Y(_130_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf2), .C(z_3_), .Y(_131_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_130_), .C(_131_), .Y(_20__3_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_4_), .Y(_132_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf0), .B(_124__bF_buf2), .C(z_4_), .Y(_133_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_132_), .C(_133_), .Y(_20__4_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_5_), .Y(_134_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_5_), .Y(_135_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_134_), .C(_135_), .Y(_20__5_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_6_), .Y(_136_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf0), .C(z_6_), .Y(_137_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_136_), .C(_137_), .Y(_20__6_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_7_), .Y(_138_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf0), .B(_124__bF_buf2), .C(z_7_), .Y(_139_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_138_), .C(_139_), .Y(_20__7_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_8_), .Y(_140_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_8_), .Y(_141_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_140_), .C(_141_), .Y(_20__8_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_9_), .Y(_142_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf2), .B(_124__bF_buf1), .C(z_9_), .Y(_143_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_142_), .C(_143_), .Y(_20__9_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_10_), .Y(_144_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf0), .C(z_10_), .Y(_145_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_144_), .C(_145_), .Y(_20__10_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf0), .B(z_m_11_), .Y(_146_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf0), .B(_124__bF_buf1), .C(z_11_), .Y(_147_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_146_), .C(_147_), .Y(_20__11_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_12_), .Y(_148_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_12_), .Y(_149_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_148_), .C(_149_), .Y(_20__12_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf1), .B(z_m_13_), .Y(_150_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf3), .B(_124__bF_buf3), .C(z_13_), .Y(_151_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf4), .B(_150_), .C(_151_), .Y(_20__13_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_14_), .Y(_152_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf0), .B(_124__bF_buf1), .C(z_14_), .Y(_153_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_152_), .C(_153_), .Y(_20__14_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_15_), .Y(_154_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf0), .C(z_15_), .Y(_155_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_154_), .C(_155_), .Y(_20__15_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_16_), .Y(_156_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf2), .B(_124__bF_buf1), .C(z_16_), .Y(_157_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_156_), .C(_157_), .Y(_20__16_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_17_), .Y(_158_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf2), .C(z_17_), .Y(_159_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_158_), .C(_159_), .Y(_20__17_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf4), .B(z_m_18_), .Y(_160_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf0), .C(z_18_), .Y(_161_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_160_), .C(_161_), .Y(_20__18_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf0), .B(z_m_19_), .Y(_162_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf0), .C(z_19_), .Y(_163_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_162_), .C(_163_), .Y(_20__19_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_20_), .Y(_164_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf0), .B(_124__bF_buf1), .C(z_20_), .Y(_165_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf2), .B(_164_), .C(_165_), .Y(_20__20_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_21_), .Y(_166_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_38__bF_buf4), .B(_124__bF_buf2), .C(z_21_), .Y(_167_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf3), .B(_166_), .C(_167_), .Y(_20__21_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(count_0_), .Y(_168_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .B(_168_), .Y(_169_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .B(count_3_), .Y(_171_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(count_4_), .B(count_5_), .C(_171_), .Y(_172_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_170_), .Y(_173_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_173_), .C(state_1_bF_buf2), .Y(_174_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(state_6_bF_buf3), .Y(_175_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_175_), .Y(_176_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_176_), .C(_174_), .Y(_8__0_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .Y(_177_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_177_), .Y(_178_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_170_), .C(state_1_bF_buf2), .Y(_179_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .Y(_180_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .B(_175_), .C(_180_), .Y(_181_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_177_), .C(_181_), .Y(_8__1_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .Y(_182_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(_182__bF_buf5), .C(count_2_), .Y(_183_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(_178_), .Y(_184_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .Y(_185_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_184_), .Y(_186_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .C(_186_), .Y(_8__2_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(_182__bF_buf5), .C(count_3_), .Y(_187_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(count_3_), .B(_187_), .S(_186_), .Y(_8__3_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(count_3_), .B(_186_), .Y(_188_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(_182__bF_buf2), .C(count_4_), .Y(_189_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(count_4_), .Y(_190_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_188_), .Y(_191_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_189_), .C(_191_), .Y(_8__4_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .B(_182__bF_buf2), .C(count_5_), .Y(_192_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(count_5_), .B(_192_), .S(_191_), .Y(_8__5_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf6), .Y(_193_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_193_), .Y(_1953_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf1), .Y(_194_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_194__bF_buf1), .Y(_1954_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(b_m_23_), .Y(_195_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_10_), .Y(_196_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .Y(_197_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_197_), .Y(_198_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_198_), .Y(_1955_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .Y(_199_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_199__bF_buf5), .Y(_1956_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf2), .Y(_200_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_200_), .Y(_201_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_201_), .Y(_1957_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(state_8_), .B(input_b_stb), .C(_2005_), .Y(_202_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_202__bF_buf6), .Y(_1958_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_203_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(z_e_8_), .Y(_204_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(z_e_0_), .Y(_205_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(z_e_1_), .Y(_206_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .Y(_207_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(z_e_5_), .Y(_208_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(z_e_4_), .Y(_209_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(z_e_6_), .Y(_211_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(z_e_7_), .B(_211_), .Y(_212_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_210_), .Y(_213_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .B(z_e_2_), .Y(_214_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_213_), .Y(_215_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_215_), .C(z_e_7_), .Y(_216_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_216_), .C(z_e_9_), .Y(_217_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(_218_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(z_e_1_), .B(_205_), .Y(_219_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_219_), .Y(_220_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_220_), .C(_213_), .Y(_221_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_218_), .Y(_222_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(state_13_), .B(_222_), .Y(_223_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_224_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_224_), .Y(_225_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_225_), .Y(_1959_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_226_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(input_a_stb), .B(_2004_), .Y(_227_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .Y(_228_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(output_z_ack), .B(_2007_), .Y(_229_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf0), .B(_229_), .C(_203_), .Y(_230_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_230_), .Y(_231_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_227_), .C(_231_), .Y(_1960_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_182__bF_buf5), .C(rst), .Y(_1961_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .B(_218_), .C(state_5_), .Y(_232_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(state_13_), .Y(_233_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_222_), .Y(_234_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf4), .Y(_235_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_232_), .C(rst), .Y(_1962_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .Y(_236_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(b_m_23_), .B(_196_), .Y(_237_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_237__bF_buf1), .Y(_238_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_238_), .C(rst), .Y(_1963_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .Y(_239_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .Y(_240_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .B(_218_), .Y(_241_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_241_), .Y(_242_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_242_), .Y(_243_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf0), .Y(_244_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_239__bF_buf2), .C(rst), .Y(_1964_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_227_), .Y(_245_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(input_b_stb), .B(_2005_), .Y(_246_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(state_8_), .B(_246_), .Y(_247_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_245__bF_buf4), .B(_247_), .C(rst), .Y(_1965_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_1974__bF_buf0), .Y(_248_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_124__bF_buf2), .Y(_249_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_248_), .C(rst), .Y(_1966_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_51_), .Y(_250_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_123_), .C(state_12_bF_buf1), .Y(_251_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(state_7_bF_buf2), .C(state_11_bF_buf0), .Y(_252_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_252_), .C(rst), .Y(_1967_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(divisor_0_), .Y(_253_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_0_), .Y(_254_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(_253_), .C(_254_), .Y(_10__0_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(divisor_1_), .Y(_255_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(b_m_1_), .Y(_256_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_255_), .C(_256_), .Y(_10__1_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(b_m_2_), .Y(_257_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(divisor_2_), .B(_182__bF_buf3), .Y(_258_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf3), .B(_257_), .C(_258_), .Y(_10__2_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(b_m_3_), .Y(_259_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(divisor_3_), .B(_182__bF_buf3), .Y(_260_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf3), .B(_259_), .C(_260_), .Y(_10__3_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(b_m_4_), .Y(_261_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(divisor_4_), .B(_182__bF_buf3), .Y(_262_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf0), .B(_261_), .C(_262_), .Y(_10__4_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(divisor_5_), .Y(_263_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(b_m_5_), .Y(_264_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(_263_), .C(_264_), .Y(_10__5_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(divisor_6_), .B(_182__bF_buf3), .Y(_265_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf3), .B(_66_), .C(_265_), .Y(_10__6_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(divisor_7_), .Y(_266_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_7_), .Y(_267_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_266_), .C(_267_), .Y(_10__7_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(divisor_8_), .Y(_268_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_8_), .Y(_269_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_268_), .C(_269_), .Y(_10__8_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(divisor_9_), .Y(_270_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(b_m_9_), .Y(_271_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_270_), .C(_271_), .Y(_10__9_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(b_m_10_), .Y(_272_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(divisor_10_), .B(_182__bF_buf2), .Y(_273_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf2), .B(_272_), .C(_273_), .Y(_10__10_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(divisor_11_), .Y(_274_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_11_), .Y(_275_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_274_), .C(_275_), .Y(_10__11_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(divisor_12_), .Y(_276_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_12_), .Y(_277_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf2), .B(_276_), .C(_277_), .Y(_10__12_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(divisor_13_), .Y(_278_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(b_m_13_), .Y(_279_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf7), .B(_278_), .C(_279_), .Y(_10__13_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(divisor_14_), .Y(_280_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_14_), .Y(_281_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(_280_), .C(_281_), .Y(_10__14_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(divisor_15_), .Y(_282_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_15_), .Y(_283_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_282_), .C(_283_), .Y(_10__15_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(divisor_16_), .Y(_284_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_16_), .Y(_285_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_284_), .C(_285_), .Y(_10__16_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(divisor_17_), .Y(_286_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_17_), .Y(_287_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_286_), .C(_287_), .Y(_10__17_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(divisor_18_), .Y(_288_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_18_), .Y(_289_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_288_), .C(_289_), .Y(_10__18_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(divisor_19_), .Y(_290_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(b_m_19_), .Y(_291_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf0), .B(_290_), .C(_291_), .Y(_10__19_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(divisor_20_), .Y(_292_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(b_m_20_), .Y(_293_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(_292_), .C(_293_), .Y(_10__20_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(divisor_21_), .Y(_294_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(b_m_21_), .Y(_295_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(_294_), .C(_295_), .Y(_10__21_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(b_m_22_), .Y(_296_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(divisor_22_), .B(_182__bF_buf2), .Y(_297_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf5), .B(_296_), .C(_297_), .Y(_10__22_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(divisor_23_), .Y(_298_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(b_m_23_), .Y(_299_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(_298_), .C(_299_), .Y(_10__23_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(divisor_24_), .Y(_300_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_300_), .Y(_10__24_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(divisor_25_), .Y(_301_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_301_), .Y(_10__25_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(divisor_26_), .Y(_302_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_302_), .Y(_10__26_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(divisor_27_), .Y(_303_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_303_), .Y(_10__27_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(divisor_28_), .Y(_304_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_304_), .Y(_10__28_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(divisor_29_), .Y(_305_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf6), .B(_305_), .Y(_10__29_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(divisor_30_), .Y(_306_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_306_), .Y(_10__30_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(divisor_31_), .Y(_307_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_307_), .Y(_10__31_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(divisor_32_), .Y(_308_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_308_), .Y(_10__32_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(divisor_33_), .Y(_309_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_309_), .Y(_10__33_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(divisor_34_), .Y(_310_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf3), .B(_310_), .Y(_10__34_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(divisor_35_), .Y(_311_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_311_), .Y(_10__35_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(divisor_36_), .Y(_312_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_312_), .Y(_10__36_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(divisor_37_), .Y(_313_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_313_), .Y(_10__37_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(divisor_38_), .Y(_314_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_314_), .Y(_10__38_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(divisor_39_), .Y(_315_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_315_), .Y(_10__39_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(divisor_40_), .Y(_316_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_316_), .Y(_10__40_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(divisor_41_), .Y(_317_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_317_), .Y(_10__41_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf2), .B(divisor_42_), .Y(_10__42_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(divisor_43_), .Y(_318_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_318_), .Y(_10__43_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf2), .B(divisor_44_), .Y(_10__44_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(divisor_45_), .Y(_319_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_319_), .Y(_10__45_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(divisor_46_), .Y(_320_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_320_), .Y(_10__46_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(divisor_47_), .Y(_321_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf1), .B(_321_), .Y(_10__47_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(divisor_48_), .Y(_322_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_322_), .Y(_10__48_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(divisor_49_), .Y(_323_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf4), .B(_323_), .Y(_10__49_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(divisor_50_), .Y(_324_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf3), .B(_324_), .Y(_10__50_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(a_s), .B(b_s), .Y(_325_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_325_), .Y(_326_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(z_s), .B(_182__bF_buf4), .Y(_327_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf4), .B(_326_), .C(_327_), .Y(_23_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(b_31_), .Y(_328_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(b_s), .B(_193_), .Y(_329_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_328_), .C(_329_), .Y(_7_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(a_31_), .Y(_330_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(a_s), .B(_193_), .Y(_331_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_330_), .C(_331_), .Y(_3_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(b_0_), .Y(_332_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(input_b[0]), .B(_202__bF_buf0), .Y(_333_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_202__bF_buf1), .C(_333_), .Y(_4__0_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(b_1_), .Y(_334_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(input_b[1]), .B(_202__bF_buf1), .Y(_335_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_202__bF_buf1), .C(_335_), .Y(_4__1_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(b_2_), .Y(_336_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(input_b[2]), .B(_202__bF_buf3), .Y(_337_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_202__bF_buf3), .C(_337_), .Y(_4__2_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(b_3_), .Y(_338_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(input_b[3]), .B(_202__bF_buf2), .Y(_339_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_202__bF_buf1), .C(_339_), .Y(_4__3_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(b_4_), .Y(_340_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(input_b[4]), .B(_202__bF_buf2), .Y(_341_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_202__bF_buf1), .C(_341_), .Y(_4__4_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(b_5_), .Y(_342_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(input_b[5]), .B(_202__bF_buf3), .Y(_343_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_202__bF_buf2), .C(_343_), .Y(_4__5_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(b_6_), .Y(_344_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(input_b[6]), .B(_202__bF_buf7), .Y(_345_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_202__bF_buf4), .C(_345_), .Y(_4__6_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(b_7_), .Y(_346_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(input_b[7]), .B(_202__bF_buf2), .Y(_347_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_202__bF_buf4), .C(_347_), .Y(_4__7_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(b_8_), .Y(_348_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(input_b[8]), .B(_202__bF_buf4), .Y(_349_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_202__bF_buf4), .C(_349_), .Y(_4__8_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(b_9_), .Y(_350_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(input_b[9]), .B(_202__bF_buf7), .Y(_351_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_202__bF_buf7), .C(_351_), .Y(_4__9_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(b_10_), .Y(_352_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(input_b[10]), .B(_202__bF_buf7), .Y(_353_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_202__bF_buf4), .C(_353_), .Y(_4__10_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(b_11_), .Y(_354_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(input_b[11]), .B(_202__bF_buf7), .Y(_355_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_202__bF_buf7), .C(_355_), .Y(_4__11_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(b_12_), .Y(_356_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(input_b[12]), .B(_202__bF_buf2), .Y(_357_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_202__bF_buf3), .C(_357_), .Y(_4__12_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(b_13_), .Y(_358_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(input_b[13]), .B(_202__bF_buf7), .Y(_359_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_202__bF_buf4), .C(_359_), .Y(_4__13_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(b_14_), .Y(_360_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(input_b[14]), .B(_202__bF_buf7), .Y(_361_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_202__bF_buf7), .C(_361_), .Y(_4__14_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(b_15_), .Y(_362_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(input_b[15]), .B(_202__bF_buf3), .Y(_363_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_202__bF_buf4), .C(_363_), .Y(_4__15_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(b_16_), .Y(_364_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(input_b[16]), .B(_202__bF_buf1), .Y(_365_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_202__bF_buf6), .C(_365_), .Y(_4__16_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(b_17_), .Y(_366_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(input_b[17]), .B(_202__bF_buf6), .Y(_367_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_202__bF_buf6), .C(_367_), .Y(_4__17_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(b_18_), .Y(_368_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(input_b[18]), .B(_202__bF_buf0), .Y(_369_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_202__bF_buf3), .C(_369_), .Y(_4__18_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(b_19_), .Y(_370_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(input_b[19]), .B(_202__bF_buf2), .Y(_371_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_202__bF_buf4), .C(_371_), .Y(_4__19_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(b_20_), .Y(_372_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(input_b[20]), .B(_202__bF_buf2), .Y(_373_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_202__bF_buf2), .C(_373_), .Y(_4__20_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(b_21_), .Y(_374_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(input_b[21]), .B(_202__bF_buf6), .Y(_375_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_202__bF_buf5), .C(_375_), .Y(_4__21_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(b_22_), .Y(_376_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(input_b[22]), .B(_202__bF_buf3), .Y(_377_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_202__bF_buf3), .C(_377_), .Y(_4__22_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(b_23_), .Y(_378_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(input_b[23]), .B(_202__bF_buf6), .Y(_379_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_202__bF_buf6), .C(_379_), .Y(_4__23_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(b_24_), .Y(_380_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(input_b[24]), .B(_202__bF_buf5), .Y(_381_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_202__bF_buf5), .C(_381_), .Y(_4__24_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(b_25_), .Y(_382_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(input_b[25]), .B(_202__bF_buf6), .Y(_383_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_202__bF_buf5), .C(_383_), .Y(_4__25_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(b_26_), .Y(_384_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(input_b[26]), .B(_202__bF_buf0), .Y(_385_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_202__bF_buf1), .C(_385_), .Y(_4__26_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(b_27_), .Y(_386_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(input_b[27]), .B(_202__bF_buf0), .Y(_387_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_202__bF_buf5), .C(_387_), .Y(_4__27_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(b_28_), .Y(_388_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(input_b[28]), .B(_202__bF_buf0), .Y(_389_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_202__bF_buf1), .C(_389_), .Y(_4__28_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(b_29_), .Y(_390_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(input_b[29]), .B(_202__bF_buf0), .Y(_391_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_202__bF_buf5), .C(_391_), .Y(_4__29_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(b_30_), .Y(_392_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(input_b[30]), .B(_202__bF_buf5), .Y(_393_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_202__bF_buf5), .C(_393_), .Y(_4__30_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(input_b[31]), .B(_202__bF_buf0), .Y(_394_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_202__bF_buf6), .C(_394_), .Y(_4__31_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(a_0_), .Y(_395_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(input_a[0]), .B(_245__bF_buf2), .Y(_396_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_245__bF_buf2), .C(_396_), .Y(_0__0_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(a_1_), .Y(_397_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(input_a[1]), .B(_245__bF_buf7), .Y(_398_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_245__bF_buf7), .C(_398_), .Y(_0__1_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(a_2_), .Y(_399_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(input_a[2]), .B(_245__bF_buf1), .Y(_400_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_245__bF_buf3), .C(_400_), .Y(_0__2_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(a_3_), .Y(_401_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(input_a[3]), .B(_245__bF_buf2), .Y(_402_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_245__bF_buf3), .C(_402_), .Y(_0__3_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(a_4_), .Y(_403_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(input_a[4]), .B(_245__bF_buf3), .Y(_404_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_245__bF_buf3), .C(_404_), .Y(_0__4_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(a_5_), .Y(_405_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(input_a[5]), .B(_245__bF_buf1), .Y(_406_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_245__bF_buf5), .C(_406_), .Y(_0__5_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(a_6_), .Y(_407_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(input_a[6]), .B(_245__bF_buf7), .Y(_408_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_245__bF_buf5), .C(_408_), .Y(_0__6_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(a_7_), .Y(_409_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(input_a[7]), .B(_245__bF_buf5), .Y(_410_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_245__bF_buf7), .C(_410_), .Y(_0__7_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(a_8_), .Y(_411_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(input_a[8]), .B(_245__bF_buf5), .Y(_412_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_245__bF_buf5), .C(_412_), .Y(_0__8_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(a_9_), .Y(_413_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(input_a[9]), .B(_245__bF_buf1), .Y(_414_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_245__bF_buf1), .C(_414_), .Y(_0__9_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(a_10_), .Y(_415_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(input_a[10]), .B(_245__bF_buf7), .Y(_416_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_245__bF_buf7), .C(_416_), .Y(_0__10_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(a_11_), .Y(_417_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(input_a[11]), .B(_245__bF_buf2), .Y(_418_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_245__bF_buf2), .C(_418_), .Y(_0__11_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(a_12_), .Y(_419_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(input_a[12]), .B(_245__bF_buf2), .Y(_420_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_245__bF_buf4), .C(_420_), .Y(_0__12_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(a_13_), .Y(_421_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(input_a[13]), .B(_245__bF_buf4), .Y(_422_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_245__bF_buf4), .C(_422_), .Y(_0__13_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(a_14_), .Y(_423_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(input_a[14]), .B(_245__bF_buf4), .Y(_424_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_245__bF_buf4), .C(_424_), .Y(_0__14_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(a_15_), .Y(_425_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(input_a[15]), .B(_245__bF_buf2), .Y(_426_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_245__bF_buf2), .C(_426_), .Y(_0__15_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(a_16_), .Y(_427_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(input_a[16]), .B(_245__bF_buf3), .Y(_428_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_245__bF_buf3), .C(_428_), .Y(_0__16_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(a_17_), .Y(_429_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(input_a[17]), .B(_245__bF_buf1), .Y(_430_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_245__bF_buf3), .C(_430_), .Y(_0__17_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(a_18_), .Y(_431_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(input_a[18]), .B(_245__bF_buf5), .Y(_432_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_245__bF_buf6), .C(_432_), .Y(_0__18_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(a_19_), .Y(_433_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(input_a[19]), .B(_245__bF_buf1), .Y(_434_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_245__bF_buf3), .C(_434_), .Y(_0__19_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(a_20_), .Y(_435_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(input_a[20]), .B(_245__bF_buf7), .Y(_436_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_245__bF_buf6), .C(_436_), .Y(_0__20_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(a_21_), .Y(_437_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(input_a[21]), .B(_245__bF_buf1), .Y(_438_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_245__bF_buf5), .C(_438_), .Y(_0__21_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(a_22_), .Y(_439_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(input_a[22]), .B(_245__bF_buf7), .Y(_440_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_245__bF_buf7), .C(_440_), .Y(_0__22_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(a_23_), .Y(_441_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(input_a[23]), .B(_245__bF_buf6), .Y(_442_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_245__bF_buf6), .C(_442_), .Y(_0__23_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(a_24_), .Y(_443_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(input_a[24]), .B(_245__bF_buf1), .Y(_444_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_245__bF_buf6), .C(_444_), .Y(_0__24_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(a_25_), .Y(_445_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(input_a[25]), .B(_245__bF_buf0), .Y(_446_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_245__bF_buf0), .C(_446_), .Y(_0__25_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(a_26_), .Y(_447_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(input_a[26]), .B(_245__bF_buf4), .Y(_448_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_245__bF_buf4), .C(_448_), .Y(_0__26_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(a_27_), .Y(_449_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(input_a[27]), .B(_245__bF_buf0), .Y(_450_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_245__bF_buf0), .C(_450_), .Y(_0__27_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(a_28_), .Y(_451_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(input_a[28]), .B(_245__bF_buf6), .Y(_452_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_245__bF_buf6), .C(_452_), .Y(_0__28_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(a_29_), .Y(_453_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(input_a[29]), .B(_245__bF_buf0), .Y(_454_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_245__bF_buf0), .C(_454_), .Y(_0__29_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(a_30_), .Y(_455_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(input_a[30]), .B(_245__bF_buf0), .Y(_456_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_245__bF_buf0), .C(_456_), .Y(_0__30_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(input_a[31]), .B(_245__bF_buf5), .Y(_457_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_245__bF_buf6), .C(_457_), .Y(_0__31_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(state_8_), .B(_2005_), .C(_202__bF_buf0), .Y(_458_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_458_), .Y(_16_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_2004_), .C(_245__bF_buf6), .Y(_459_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_459_), .Y(_15_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_2006__0_), .Y(_460_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(z_0_), .B(state_7_bF_buf5), .Y(_461_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_460_), .C(_461_), .Y(_17__0_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(_2006__1_), .Y(_462_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(z_1_), .B(state_7_bF_buf0), .Y(_463_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf3), .B(_462_), .C(_463_), .Y(_17__1_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_2006__2_), .Y(_464_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(z_2_), .B(state_7_bF_buf4), .Y(_465_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf4), .B(_464_), .C(_465_), .Y(_17__2_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_2006__3_), .Y(_466_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(z_3_), .B(state_7_bF_buf0), .Y(_467_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf2), .B(_466_), .C(_467_), .Y(_17__3_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_2006__4_), .Y(_468_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(z_4_), .B(state_7_bF_buf0), .Y(_469_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf2), .B(_468_), .C(_469_), .Y(_17__4_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_2006__5_), .Y(_470_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(z_5_), .B(state_7_bF_buf0), .Y(_471_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf5), .B(_470_), .C(_471_), .Y(_17__5_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_2006__6_), .Y(_472_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(z_6_), .B(state_7_bF_buf3), .Y(_473_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf3), .B(_472_), .C(_473_), .Y(_17__6_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_2006__7_), .Y(_474_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(z_7_), .B(state_7_bF_buf0), .Y(_475_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_474_), .C(_475_), .Y(_17__7_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_2006__8_), .Y(_476_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(z_8_), .B(state_7_bF_buf3), .Y(_477_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf5), .B(_476_), .C(_477_), .Y(_17__8_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_2006__9_), .Y(_478_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(z_9_), .B(state_7_bF_buf4), .Y(_479_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf4), .B(_478_), .C(_479_), .Y(_17__9_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_2006__10_), .Y(_480_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(z_10_), .B(state_7_bF_buf3), .Y(_481_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_480_), .C(_481_), .Y(_17__10_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_2006__11_), .Y(_482_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(z_11_), .B(state_7_bF_buf2), .Y(_483_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_482_), .C(_483_), .Y(_17__11_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_2006__12_), .Y(_484_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(z_12_), .B(state_7_bF_buf3), .Y(_485_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_484_), .C(_485_), .Y(_17__12_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_2006__13_), .Y(_486_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(z_13_), .B(state_7_bF_buf3), .Y(_487_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_486_), .C(_487_), .Y(_17__13_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_2006__14_), .Y(_488_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(z_14_), .B(state_7_bF_buf2), .Y(_489_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf4), .B(_488_), .C(_489_), .Y(_17__14_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_2006__15_), .Y(_490_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(z_15_), .B(state_7_bF_buf5), .Y(_491_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf5), .B(_490_), .C(_491_), .Y(_17__15_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_2006__16_), .Y(_492_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(z_16_), .B(state_7_bF_buf4), .Y(_493_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf4), .B(_492_), .C(_493_), .Y(_17__16_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_2006__17_), .Y(_494_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(z_17_), .B(state_7_bF_buf0), .Y(_495_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_494_), .C(_495_), .Y(_17__17_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_2006__18_), .Y(_496_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(z_18_), .B(state_7_bF_buf5), .Y(_497_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_496_), .C(_497_), .Y(_17__18_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_2006__19_), .Y(_498_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(z_19_), .B(state_7_bF_buf6), .Y(_499_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf6), .B(_498_), .C(_499_), .Y(_17__19_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_2006__20_), .Y(_500_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(z_20_), .B(state_7_bF_buf2), .Y(_501_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf2), .B(_500_), .C(_501_), .Y(_17__20_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_2006__21_), .Y(_502_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(z_21_), .B(state_7_bF_buf0), .Y(_503_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf5), .B(_502_), .C(_503_), .Y(_17__21_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_2006__22_), .Y(_504_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(z_22_), .Y(_505_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_504_), .C(_505_), .Y(_17__22_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(z_23_), .Y(_506_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_2006__23_), .B(_228__bF_buf3), .Y(_507_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf3), .B(_506_), .C(_507_), .Y(_17__23_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(z_24_), .Y(_508_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_2006__24_), .B(_228__bF_buf0), .Y(_509_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf2), .B(_508_), .C(_509_), .Y(_17__24_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(z_25_), .Y(_510_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_2006__25_), .B(_228__bF_buf0), .Y(_511_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf2), .B(_510_), .C(_511_), .Y(_17__25_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(z_26_), .Y(_512_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_2006__26_), .B(_228__bF_buf3), .Y(_513_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf3), .B(_512_), .C(_513_), .Y(_17__26_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(z_27_), .Y(_514_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2006__27_), .B(_228__bF_buf1), .Y(_515_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf1), .B(_514_), .C(_515_), .Y(_17__27_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(z_28_), .Y(_516_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_2006__28_), .B(_228__bF_buf2), .Y(_517_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf2), .B(_516_), .C(_517_), .Y(_17__28_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(z_29_), .Y(_518_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_2006__29_), .B(_228__bF_buf1), .Y(_519_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf1), .B(_518_), .C(_519_), .Y(_17__29_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(z_30_), .Y(_520_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_2006__30_), .B(_228__bF_buf0), .Y(_521_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf3), .B(_520_), .C(_521_), .Y(_17__30_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_2006__31_), .Y(_522_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(z_31_), .Y(_523_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_522_), .C(_523_), .Y(_17__31_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .Y(_524_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_228__bF_buf2), .B(_524_), .C(_230_), .Y(_18_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_86_), .Y(_525_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_109_), .Y(_526_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_118_), .Y(_527_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_527_), .Y(_528_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_528_), .Y(_529_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_526_), .Y(_530_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_525_), .Y(_531_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_528_), .Y(_532_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_532_), .Y(_533_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_533_), .Y(_534_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_91_), .Y(_535_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(_535_), .Y(_536_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_51_), .C(z_22_), .Y(_537_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_536_), .C(_122_), .Y(_538_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_537_), .C(_538_), .Y(_539_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_539_), .C(state_12_bF_buf2), .Y(_540_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(z_22_), .B(_38__bF_buf0), .Y(_541_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf3), .B(z_m_22_), .C(_35_), .Y(_542_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_542_), .C(_540_), .Y(_20__22_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(z_m_0_), .Y(_543_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(state_13_), .B(state_5_), .Y(_544_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf2), .B(_544_), .Y(_545_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_223_), .Y(_546_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_546_), .Y(_547_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf1), .B(_545_), .C(_547_), .Y(_548_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_548_), .Y(_549_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(z_m_1_), .B(_234__bF_buf1), .Y(_550_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(quotient_3_), .Y(_551_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(guard), .Y(_552_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(round_bit), .B(sticky), .Y(_553_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_543_), .C(_552_), .Y(_554_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(z_m_0_), .B(guard), .C(_194__bF_buf3), .Y(_555_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(z_m_0_), .B(_554_), .C(_555_), .Y(_556_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf3), .B(_551_), .C(_556_), .Y(_557_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf2), .B(guard), .C(_557_), .Y(_558_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_550_), .Y(_559_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_549_), .C(_559_), .Y(_22__0_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(quotient_0_), .Y(_560_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(state_14_bF_buf7), .Y(_561_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(_561__bF_buf4), .Y(_562_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(state_1_bF_buf1), .B(_562__bF_buf4), .Y(_563_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_563__bF_buf2), .Y(_564_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(remainder_50_), .Y(_565_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(divisor_50_), .B(_565_), .Y(_566_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_566_), .Y(_567_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(remainder_46_), .B(_320_), .Y(_568_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(remainder_46_), .B(_320_), .Y(_569_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_569_), .Y(_570_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_570_), .Y(_571_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(remainder_47_), .Y(_572_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(divisor_47_), .B(_572_), .Y(_573_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(remainder_47_), .B(_321_), .Y(_574_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_574_), .Y(_575_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_571_), .Y(_576_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(remainder_45_), .Y(_577_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(remainder_45_), .B(_319_), .Y(_578_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_577_), .Y(_579_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(remainder_44_), .Y(_580_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(divisor_44_), .B(_580_), .Y(_581_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_581_), .Y(_582_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(divisor_44_), .B(_580_), .Y(_583_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_582_), .Y(_584_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_584_), .Y(_585_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_585_), .Y(_586_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_586_), .Y(_587_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(remainder_42_), .Y(_588_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(divisor_42_), .B(_588_), .Y(_589_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(divisor_42_), .B(_588_), .Y(_590_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_590_), .Y(_591_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(remainder_43_), .Y(_592_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(divisor_43_), .B(_592_), .Y(_593_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(remainder_43_), .B(_318_), .Y(_594_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_594_), .Y(_595_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_591_), .C(_595_), .Y(_596_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(remainder_41_), .Y(_597_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(divisor_41_), .B(_597_), .Y(_598_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_598_), .Y(_599_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(remainder_40_), .B(_316_), .Y(_600_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(remainder_41_), .B(_317_), .Y(_601_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_601_), .C(_599_), .Y(_602_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_602_), .Y(_603_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_590_), .C(_593_), .Y(_604_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_603_), .C(_604_), .Y(_605_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_581_), .C(_577_), .Y(_606_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_570_), .C(_573_), .Y(_607_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_606_), .C(_607_), .Y(_608_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_587_), .C(_608_), .Y(_609_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_601_), .Y(_610_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_610_), .Y(_611_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(remainder_40_), .Y(_612_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(divisor_40_), .B(_612_), .Y(_613_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_613_), .Y(_614_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_614_), .Y(_615_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_611_), .Y(_616_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_616_), .Y(_617_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_617_), .Y(_618_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_587_), .Y(_619_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(divisor_38_), .B(remainder_38_), .Y(_620_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(remainder_39_), .Y(_621_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(divisor_39_), .B(_621_), .Y(_622_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(remainder_39_), .B(_315_), .Y(_623_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_623_), .Y(_624_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_624_), .Y(_625_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_625_), .Y(_626_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(remainder_37_), .Y(_627_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(remainder_36_), .B(_312_), .Y(_628_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(divisor_37_), .B(_627_), .C(_628_), .Y(_629_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(remainder_37_), .C(_629_), .Y(_630_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_630_), .Y(_631_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_620_), .Y(_632_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(remainder_37_), .B(_313_), .Y(_633_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(divisor_37_), .B(_627_), .Y(_634_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_634_), .Y(_635_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(remainder_36_), .Y(_636_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(divisor_36_), .B(_636_), .Y(_637_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_637_), .Y(_638_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_635_), .Y(_639_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_624_), .C(_639_), .Y(_640_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(remainder_34_), .Y(_641_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(remainder_34_), .B(_310_), .Y(_642_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_641_), .Y(_643_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(remainder_35_), .Y(_644_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(divisor_35_), .B(_644_), .Y(_645_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(remainder_35_), .B(_311_), .Y(_646_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_646_), .Y(_647_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_648_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_648_), .Y(_649_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(remainder_33_), .B(_309_), .Y(_650_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(remainder_32_), .B(_308_), .Y(_651_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(remainder_33_), .Y(_652_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(divisor_33_), .B(_652_), .Y(_653_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_650_), .Y(_654_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_654_), .C(_650_), .Y(_655_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_642_), .Y(_656_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(remainder_35_), .C(_656_), .Y(_657_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(divisor_35_), .B(_644_), .C(_657_), .Y(_658_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_655_), .C(_658_), .Y(_659_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(remainder_38_), .B(_314_), .Y(_660_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(divisor_39_), .B(_621_), .C(_660_), .Y(_661_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(remainder_39_), .C(_661_), .Y(_662_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_659_), .C(_662_), .Y(_663_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_631_), .C(_663_), .Y(_664_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(remainder_1_), .B(_255_), .Y(_665_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(_665_), .Y(_666_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(remainder_0_), .Y(_667_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(remainder_1_), .Y(_668_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(divisor_1_), .B(_668_), .Y(_669_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_669_), .C(_666_), .Y(_670_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(remainder_3_), .Y(_671_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(divisor_3_), .B(_671_), .Y(_672_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(remainder_2_), .Y(_673_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(divisor_2_), .B(_673_), .Y(_674_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(divisor_3_), .B(remainder_3_), .Y(_675_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_674_), .C(_672_), .Y(_676_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(divisor_2_), .B(remainder_2_), .Y(_677_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_675_), .Y(_678_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_670_), .C(_676_), .Y(_679_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(remainder_7_), .Y(_680_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(divisor_7_), .B(_680_), .Y(_681_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(remainder_6_), .Y(_682_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(divisor_6_), .B(_682_), .Y(_683_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(divisor_7_), .B(remainder_7_), .Y(_684_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_680_), .Y(_685_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_685_), .Y(_686_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_683_), .C(_681_), .Y(_687_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(divisor_6_), .B(remainder_6_), .Y(_688_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_686_), .Y(_689_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(remainder_5_), .Y(_690_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(divisor_5_), .B(_690_), .Y(_691_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(remainder_4_), .Y(_692_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(divisor_4_), .B(_692_), .Y(_693_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(divisor_5_), .B(remainder_5_), .Y(_694_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_693_), .C(_691_), .Y(_695_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_695_), .C(_687_), .Y(_696_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(divisor_6_), .B(remainder_6_), .Y(_697_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_685_), .C(_697_), .Y(_698_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(divisor_5_), .B(remainder_5_), .Y(_699_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(divisor_4_), .B(remainder_4_), .Y(_700_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_700_), .Y(_701_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_698_), .Y(_702_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_679_), .C(_696_), .Y(_703_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(remainder_15_), .B(_282_), .Y(_704_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(remainder_15_), .Y(_705_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(divisor_15_), .B(_705_), .Y(_706_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_706_), .Y(_707_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(divisor_14_), .B(remainder_14_), .Y(_708_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_707_), .Y(_709_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(remainder_12_), .B(_276_), .Y(_710_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(remainder_12_), .Y(_711_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(divisor_12_), .B(_711_), .Y(_712_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_712_), .Y(_713_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(remainder_13_), .B(_278_), .Y(_714_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(remainder_13_), .Y(_715_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(divisor_13_), .B(_715_), .Y(_716_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_716_), .Y(_717_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_717_), .Y(_718_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_718_), .Y(_719_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(remainder_11_), .B(_274_), .Y(_720_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(remainder_11_), .Y(_721_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(divisor_11_), .B(_721_), .Y(_722_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_722_), .Y(_723_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(divisor_10_), .B(remainder_10_), .Y(_724_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_723_), .Y(_725_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(remainder_8_), .B(_268_), .Y(_726_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(remainder_8_), .Y(_727_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(divisor_8_), .B(_727_), .Y(_728_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_728_), .Y(_729_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(divisor_9_), .B(remainder_9_), .Y(_730_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_729_), .Y(_731_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_731_), .Y(_732_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_732_), .Y(_733_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_709_), .Y(_734_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(divisor_10_), .B(remainder_10_), .Y(_735_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_722_), .C(_735_), .Y(_736_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(remainder_9_), .Y(_737_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(divisor_9_), .B(_737_), .C(_726_), .Y(_738_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(remainder_9_), .C(_738_), .Y(_739_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(remainder_10_), .Y(_740_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(divisor_10_), .B(_740_), .Y(_741_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(remainder_11_), .C(_741_), .Y(_742_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_720_), .Y(_743_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_736_), .C(_743_), .Y(_744_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_708_), .Y(_745_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(divisor_13_), .B(_715_), .C(_710_), .Y(_746_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(remainder_13_), .C(_746_), .Y(_747_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_704_), .Y(_748_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(remainder_14_), .Y(_749_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_748_), .C(_706_), .Y(_750_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_745_), .C(_750_), .Y(_751_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_744_), .C(_751_), .Y(_752_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_703_), .C(_752_), .Y(_753_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(remainder_31_), .B(_307_), .Y(_754_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(remainder_31_), .Y(_755_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(divisor_31_), .B(_755_), .Y(_756_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_756_), .Y(_757_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(divisor_30_), .B(remainder_30_), .Y(_758_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_757_), .Y(_759_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(divisor_29_), .B(remainder_29_), .Y(_760_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(remainder_28_), .B(_304_), .Y(_761_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(remainder_28_), .Y(_762_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(divisor_28_), .B(_762_), .Y(_763_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_763_), .Y(_764_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_764_), .Y(_765_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_759_), .Y(_766_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(divisor_25_), .B(remainder_25_), .Y(_767_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(remainder_24_), .B(_300_), .Y(_768_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(remainder_24_), .Y(_769_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(divisor_24_), .B(_769_), .Y(_770_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_770_), .Y(_771_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_767_), .Y(_772_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(divisor_27_), .B(remainder_27_), .Y(_773_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(divisor_26_), .B(remainder_26_), .Y(_774_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_774_), .Y(_775_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_772_), .Y(_776_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_776_), .Y(_777_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(remainder_23_), .B(_298_), .Y(_778_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(remainder_23_), .Y(_779_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(divisor_23_), .B(_779_), .Y(_780_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(divisor_22_), .B(remainder_22_), .Y(_781_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_780_), .C(_781_), .Y(_782_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(divisor_21_), .B(remainder_21_), .Y(_783_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(remainder_20_), .B(_292_), .Y(_784_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(remainder_20_), .Y(_785_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(divisor_20_), .B(_785_), .Y(_786_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_786_), .Y(_787_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_783_), .Y(_788_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_788_), .Y(_789_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(remainder_19_), .B(_290_), .Y(_790_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(remainder_19_), .Y(_791_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(divisor_19_), .B(_791_), .Y(_792_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_792_), .Y(_793_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(remainder_18_), .B(_288_), .Y(_794_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(remainder_18_), .Y(_795_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(divisor_18_), .B(_795_), .Y(_796_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_796_), .Y(_797_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_793_), .Y(_798_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(remainder_17_), .B(_286_), .Y(_799_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(remainder_17_), .Y(_800_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(divisor_17_), .B(_800_), .Y(_801_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_801_), .Y(_802_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(remainder_16_), .B(_284_), .Y(_803_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(remainder_16_), .Y(_804_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(divisor_16_), .B(_804_), .Y(_805_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_803_), .B(_805_), .Y(_806_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_802_), .Y(_807_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_807_), .Y(_808_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_789_), .Y(_809_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_809_), .Y(_810_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_792_), .Y(_811_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_796_), .Y(_812_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_811_), .Y(_813_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(divisor_19_), .B(_791_), .C(_794_), .Y(_814_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(remainder_19_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(divisor_17_), .B(_800_), .C(_803_), .Y(_816_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(remainder_17_), .C(_816_), .Y(_817_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_813_), .C(_815_), .Y(_818_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(remainder_21_), .Y(_819_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(divisor_21_), .B(_819_), .C(_784_), .Y(_820_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(remainder_21_), .C(_820_), .Y(_821_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(remainder_22_), .Y(_822_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(divisor_22_), .B(_822_), .Y(_823_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(remainder_23_), .C(_823_), .Y(_824_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_778_), .Y(_825_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_782_), .C(_825_), .Y(_826_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_789_), .C(_826_), .Y(_827_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(remainder_25_), .Y(_828_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(divisor_25_), .B(_828_), .C(_768_), .Y(_829_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(remainder_25_), .C(_829_), .Y(_830_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(remainder_27_), .Y(_831_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(remainder_26_), .Y(_832_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(divisor_26_), .B(_832_), .C(divisor_27_), .D(_831_), .Y(_833_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(remainder_27_), .C(_833_), .Y(_834_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_830_), .C(_834_), .Y(_835_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(remainder_30_), .Y(_836_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(remainder_31_), .C(_836_), .Y(_837_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(remainder_29_), .B(_305_), .Y(_838_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(remainder_29_), .B(_305_), .Y(_839_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_839_), .C(_838_), .Y(_840_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_759_), .Y(_841_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_837_), .C(_841_), .Y(_842_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_835_), .C(_842_), .Y(_843_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_827_), .C(_843_), .Y(_844_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_810_), .C(_844_), .Y(_845_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(remainder_32_), .Y(_846_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(divisor_32_), .B(_846_), .Y(_847_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_847_), .Y(_848_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_654_), .Y(_849_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_649_), .Y(_850_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_850_), .Y(_851_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_851_), .Y(_852_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_845_), .C(_664_), .Y(_853_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_853_), .Y(_854_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_854_), .Y(_855_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(remainder_49_), .Y(_856_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(divisor_49_), .B(_856_), .Y(_857_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_857_), .Y(_858_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(remainder_49_), .B(_323_), .Y(_859_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(remainder_48_), .B(_322_), .Y(_860_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_859_), .C(_858_), .Y(_861_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(remainder_48_), .Y(_862_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(divisor_48_), .B(_862_), .Y(_863_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_863_), .Y(_864_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_864_), .Y(_865_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_859_), .Y(_866_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_866_), .Y(_867_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_867_), .Y(_868_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_868_), .C(_861_), .Y(_869_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(remainder_50_), .B(_324_), .Y(_870_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_870_), .B(_869_), .C(_567__bF_buf2), .Y(_871_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(quotient_0_), .B(_871__bF_buf0), .C(state_1_bF_buf1), .Y(_872_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_564_), .C(_872_), .Y(_12__0_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(quotient_1_), .Y(_873_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_560_), .C(_873_), .D(_562__bF_buf4), .Y(_12__1_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(quotient_2_), .Y(_874_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_873_), .C(_874_), .D(_562__bF_buf4), .Y(_12__2_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_874_), .C(_551_), .D(_562__bF_buf1), .Y(_12__3_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(quotient_4_), .Y(_875_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_551_), .C(_875_), .D(_562__bF_buf1), .Y(_12__4_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(quotient_5_), .Y(_876_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_875_), .C(_876_), .D(_562__bF_buf1), .Y(_12__5_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(quotient_6_), .Y(_877_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_876_), .C(_877_), .D(_562__bF_buf1), .Y(_12__6_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(quotient_7_), .Y(_878_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_877_), .C(_878_), .D(_562__bF_buf4), .Y(_12__7_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(quotient_8_), .Y(_879_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_878_), .C(_879_), .D(_562__bF_buf4), .Y(_12__8_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(quotient_9_), .Y(_880_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_879_), .C(_880_), .D(_562__bF_buf4), .Y(_12__9_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(quotient_10_), .Y(_881_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_880_), .C(_881_), .D(_562__bF_buf4), .Y(_12__10_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(quotient_11_), .Y(_882_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_881_), .C(_882_), .D(_562__bF_buf0), .Y(_12__11_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(quotient_12_), .Y(_883_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_882_), .C(_883_), .D(_562__bF_buf0), .Y(_12__12_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(quotient_13_), .Y(_884_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_883_), .C(_884_), .D(_562__bF_buf3), .Y(_12__13_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(quotient_14_), .Y(_885_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_884_), .C(_885_), .D(_562__bF_buf2), .Y(_12__14_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(quotient_15_), .Y(_886_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_885_), .C(_886_), .D(_562__bF_buf2), .Y(_12__15_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(quotient_16_), .Y(_887_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_886_), .C(_887_), .D(_562__bF_buf2), .Y(_12__16_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(quotient_17_), .Y(_888_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_887_), .C(_888_), .D(_562__bF_buf2), .Y(_12__17_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(quotient_18_), .Y(_889_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_888_), .C(_889_), .D(_562__bF_buf2), .Y(_12__18_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(quotient_19_), .Y(_890_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_889_), .C(_890_), .D(_562__bF_buf2), .Y(_12__19_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(quotient_20_), .Y(_891_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_890_), .C(_891_), .D(_562__bF_buf0), .Y(_12__20_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(quotient_21_), .Y(_892_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_891_), .C(_892_), .D(_562__bF_buf0), .Y(_12__21_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(quotient_22_), .Y(_893_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_892_), .C(_893_), .D(_562__bF_buf0), .Y(_12__22_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(quotient_23_), .Y(_894_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_893_), .C(_894_), .D(_562__bF_buf0), .Y(_12__23_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(quotient_24_), .Y(_895_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf2), .B(_894_), .C(_895_), .D(_562__bF_buf0), .Y(_12__24_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(quotient_25_), .Y(_896_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf6), .B(_895_), .C(_896_), .D(_562__bF_buf2), .Y(_12__25_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(quotient_26_), .B(_561__bF_buf4), .Y(_897_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_896_), .C(_897_), .Y(_12__26_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_91_), .Y(_898_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf3), .Y(_899_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_4_bF_buf2), .C(_899_), .Y(_900_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(state_2_), .C(a_m_23_), .D(_900_), .Y(_901_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_80_), .C(_901_), .Y(_2__23_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf6), .B(state_10_), .Y(_902_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_197_), .Y(_903_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_332_), .C(_62_), .D(_903__bF_buf0), .Y(_6__0_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_1_), .C(b_m_0_), .D(_237__bF_buf0), .Y(_904_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_903__bF_buf0), .C(_904_), .Y(_6__1_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_2_), .C(b_m_1_), .D(_237__bF_buf2), .Y(_905_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_903__bF_buf3), .C(_905_), .Y(_6__2_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_3_), .C(b_m_2_), .D(_237__bF_buf0), .Y(_906_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_903__bF_buf0), .C(_906_), .Y(_6__3_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_4_), .C(b_m_3_), .D(_237__bF_buf0), .Y(_907_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_903__bF_buf0), .C(_907_), .Y(_6__4_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(b_m_5_), .Y(_908_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_5_), .C(b_m_4_), .D(_237__bF_buf0), .Y(_909_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_908_), .B(_903__bF_buf0), .C(_909_), .Y(_6__5_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_6_), .C(b_m_5_), .D(_237__bF_buf2), .Y(_910_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_903__bF_buf3), .C(_910_), .Y(_6__6_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_7_), .C(b_m_6_), .D(_237__bF_buf2), .Y(_911_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_903__bF_buf3), .C(_911_), .Y(_6__7_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_8_), .C(b_m_7_), .D(_237__bF_buf3), .Y(_912_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_903__bF_buf3), .C(_912_), .Y(_6__8_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_9_), .C(b_m_8_), .D(_237__bF_buf2), .Y(_913_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_903__bF_buf3), .C(_913_), .Y(_6__9_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_10_), .C(b_m_9_), .D(_237__bF_buf2), .Y(_914_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_903__bF_buf1), .C(_914_), .Y(_6__10_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(b_m_11_), .Y(_915_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf5), .B(b_11_), .C(b_m_10_), .D(_237__bF_buf2), .Y(_916_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(_903__bF_buf3), .C(_916_), .Y(_6__11_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(b_m_12_), .Y(_917_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_12_), .C(b_m_11_), .D(_237__bF_buf3), .Y(_918_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_903__bF_buf1), .C(_918_), .Y(_6__12_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(b_m_13_), .Y(_919_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_13_), .C(b_m_12_), .D(_237__bF_buf3), .Y(_920_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_903__bF_buf1), .C(_920_), .Y(_6__13_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_14_), .C(b_m_13_), .D(_237__bF_buf3), .Y(_921_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_903__bF_buf1), .C(_921_), .Y(_6__14_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_15_), .C(b_m_14_), .D(_237__bF_buf3), .Y(_922_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_903__bF_buf1), .C(_922_), .Y(_6__15_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_16_), .C(b_m_15_), .D(_237__bF_buf0), .Y(_923_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_903__bF_buf2), .C(_923_), .Y(_6__16_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_17_), .C(b_m_16_), .D(_237__bF_buf1), .Y(_924_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_903__bF_buf2), .C(_924_), .Y(_6__17_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(b_m_18_), .Y(_925_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_18_), .C(b_m_17_), .D(_237__bF_buf1), .Y(_926_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_903__bF_buf2), .C(_926_), .Y(_6__18_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(b_m_19_), .Y(_927_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf0), .B(b_19_), .C(b_m_18_), .D(_237__bF_buf3), .Y(_928_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_903__bF_buf1), .C(_928_), .Y(_6__19_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_20_), .C(b_m_19_), .D(_237__bF_buf1), .Y(_929_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_903__bF_buf2), .C(_929_), .Y(_6__20_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_21_), .C(b_m_20_), .D(_237__bF_buf1), .Y(_930_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_903__bF_buf2), .C(_930_), .Y(_6__21_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(b_22_), .C(b_m_21_), .D(_237__bF_buf1), .Y(_931_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_903__bF_buf2), .C(_931_), .Y(_6__22_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(z_m_1_), .Y(_932_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_552_), .C(_932_), .Y(_933_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_932_), .Y(_934_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(guard), .C(_194__bF_buf3), .Y(_935_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_4_), .C(_933_), .D(_935_), .Y(_936_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_244_), .C(_936_), .Y(_937_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(z_m_2_), .B(_234__bF_buf1), .C(_937_), .Y(_938_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_549_), .C(_938_), .Y(_22__1_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(z_m_2_), .Y(_939_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(_934_), .Y(_940_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_940_), .C(z_m_2_), .Y(_941_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(guard), .B(_939_), .C(_934_), .Y(_942_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_941_), .Y(_943_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_5_), .C(state_3_bF_buf4), .D(_943_), .Y(_944_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_244_), .C(_944_), .Y(_945_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(z_m_3_), .B(_234__bF_buf1), .C(_945_), .Y(_946_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_549_), .C(_946_), .Y(_22__2_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(z_m_3_), .Y(_947_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(z_m_4_), .B(_234__bF_buf1), .Y(_948_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(z_m_2_), .B(_934_), .Y(_949_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(_949_), .Y(_950_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(z_m_3_), .B(_554_), .C(_950_), .Y(_951_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_554_), .Y(_952_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_952_), .C(_947_), .Y(_953_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf4), .B(_953_), .C(_951_), .Y(_954_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf3), .B(_877_), .C(_954_), .Y(_955_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf2), .B(z_m_2_), .C(_955_), .Y(_956_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_948_), .Y(_957_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_549_), .C(_957_), .Y(_22__3_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(z_m_4_), .Y(_958_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(z_m_5_), .Y(_959_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_951_), .C(state_3_bF_buf4), .Y(_960_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_951_), .C(_960_), .Y(_961_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_7_), .C(_961_), .Y(_962_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_235_), .C(_962_), .Y(_963_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(z_m_3_), .B(_243__bF_buf2), .C(_963_), .Y(_964_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_549_), .C(_964_), .Y(_22__4_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_958_), .Y(_965_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_965_), .Y(_966_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_966_), .Y(_967_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(z_m_5_), .Y(_968_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf4), .B(_968_), .Y(_969_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf3), .B(_879_), .C(_969_), .Y(_970_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(z_m_6_), .Y(_971_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_235_), .C(_958_), .D(_244_), .Y(_972_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_972_), .Y(_973_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_549_), .C(_973_), .Y(_22__5_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(z_m_5_), .B(_966_), .Y(_974_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_974_), .C(_971_), .Y(_975_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_952_), .Y(_976_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_976_), .Y(_977_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf3), .B(_977_), .Y(_978_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_9_), .C(_975_), .D(_978_), .Y(_979_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_244_), .C(_979_), .Y(_980_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(z_m_7_), .B(_234__bF_buf2), .C(_980_), .Y(_981_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_549_), .C(_981_), .Y(_22__6_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(z_m_7_), .Y(_982_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(z_m_8_), .B(_234__bF_buf0), .Y(_983_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(z_m_7_), .C(_194__bF_buf3), .Y(_984_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(z_m_7_), .B(_977_), .C(_984_), .Y(_985_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf3), .B(_881_), .C(_985_), .Y(_986_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(z_m_6_), .B(_243__bF_buf2), .C(_986_), .Y(_987_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_983_), .Y(_988_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_549_), .C(_988_), .Y(_22__7_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(z_m_8_), .Y(_989_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(z_m_7_), .B(_977_), .Y(_990_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_989_), .Y(_991_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf3), .B(_882_), .C(_194__bF_buf3), .D(_991_), .Y(_992_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(z_m_9_), .Y(_993_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_235_), .C(_982_), .D(_244_), .Y(_994_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_992_), .Y(_995_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_549_), .C(_995_), .Y(_22__8_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(z_m_8_), .B(_243__bF_buf1), .Y(_996_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(z_m_6_), .B(z_m_7_), .C(z_m_8_), .Y(_997_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_949_), .Y(_998_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(z_m_5_), .B(_965_), .C(_998_), .Y(_999_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_999_), .Y(_1000_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(z_m_9_), .C(_194__bF_buf1), .Y(_1001_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(z_m_9_), .B(_1000_), .C(_1001_), .Y(_1002_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf0), .B(_883_), .C(_1002_), .Y(_1003_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(z_m_10_), .B(_234__bF_buf2), .C(_1003_), .Y(_1004_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_1004_), .Y(_1005_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_549_), .C(_1005_), .Y(_22__9_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(z_m_10_), .Y(_1006_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(z_m_9_), .B(_243__bF_buf1), .Y(_1007_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1008_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_1008_), .C(_1006_), .Y(_1009_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_1006_), .Y(_1010_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1000_), .Y(_1011_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf4), .B(_1011_), .C(_1009_), .Y(_1012_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf0), .B(_884_), .C(_1012_), .Y(_1013_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(z_m_11_), .B(_234__bF_buf2), .C(_1013_), .Y(_1014_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1007_), .Y(_1015_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_549_), .C(_1015_), .Y(_22__10_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(z_m_11_), .Y(_1016_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_1011_), .C(state_3_bF_buf2), .Y(_1017_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_1011_), .C(_1017_), .Y(_1018_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_14_), .C(_1018_), .Y(_1019_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(z_m_12_), .B(_234__bF_buf2), .C(z_m_10_), .D(_243__bF_buf1), .Y(_1020_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1019_), .Y(_1021_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_549_), .C(_1021_), .Y(_22__11_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_974_), .Y(_1022_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(z_m_11_), .B(_1010_), .C(_1022_), .Y(_1023_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_1023_), .Y(_1024_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(z_m_12_), .Y(_1025_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf1), .B(_545_), .Y(_1026_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .Y(_1027_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1016_), .Y(_1028_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1028_), .C(state_3_bF_buf2), .Y(_1029_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1027_), .C(_1029_), .Y(_1030_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(z_m_12_), .B(_1024_), .C(_1030_), .Y(_1031_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_15_), .C(z_m_13_), .D(_234__bF_buf2), .Y(_1032_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_244_), .C(_1032_), .Y(_1033_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(z_m_12_), .B(_546_), .C(_1033_), .Y(_1034_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1034_), .Y(_22__12_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(z_m_13_), .Y(_1035_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1028_), .C(_1035_), .Y(_1036_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1035_), .Y(_1037_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .Y(_1038_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_1028_), .Y(_1039_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .Y(_1040_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf2), .B(_1036_), .C(_1040_), .Y(_1041_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf0), .B(_887_), .C(_1025_), .D(_244_), .Y(_1042_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(z_m_14_), .B(_234__bF_buf2), .C(_1042_), .Y(_1043_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_1041_), .Y(_1044_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_549_), .C(_1044_), .Y(_22__13_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(z_m_14_), .B(_1039_), .Y(_1045_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(z_m_14_), .B(_1039_), .Y(_1046_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf2), .B(_1046_), .C(z_m_14_), .D(_548_), .Y(_1047_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(z_m_15_), .Y(_1048_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf1), .B(_888_), .C(_1048_), .D(_235_), .Y(_1049_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(z_m_13_), .B(_243__bF_buf1), .C(_1049_), .Y(_1050_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1047_), .C(_1050_), .Y(_22__14_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .Y(_1051_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_1046_), .Y(_1052_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf1), .B(_1052_), .Y(_1053_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(z_m_15_), .B(_1051_), .C(_1053_), .Y(_1054_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_546_), .C(z_m_15_), .Y(_1055_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(z_m_14_), .Y(_1056_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf0), .B(_889_), .C(_1056_), .D(_244_), .Y(_1057_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(z_m_16_), .B(_234__bF_buf0), .C(_1057_), .Y(_1058_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1058_), .C(_1054_), .Y(_22__15_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_1053_), .C(z_m_16_), .Y(_1059_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(z_m_16_), .Y(_1060_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf2), .B(_1060_), .C(_1052_), .Y(_1061_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf1), .B(_890_), .C(_1048_), .D(_244_), .Y(_1062_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(z_m_17_), .B(_234__bF_buf0), .C(_1062_), .Y(_1063_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1063_), .C(_1059_), .Y(_22__16_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_952_), .Y(_1064_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(z_m_14_), .B(_1037_), .Y(_1065_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_1065_), .Y(_1066_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(z_m_16_), .B(_1066_), .Y(_1067_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(_1064_), .Y(_1068_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(z_m_17_), .B(_1068_), .Y(_1069_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(z_m_17_), .Y(_1070_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf0), .B(_1070_), .Y(_1071_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(z_m_17_), .B(_548_), .C(_1071_), .Y(_1072_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf1), .B(_891_), .C(_1060_), .D(_244_), .Y(_1073_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(z_m_18_), .B(_234__bF_buf4), .C(_1073_), .Y(_1074_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1072_), .C(_1074_), .Y(_22__17_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_1071_), .C(z_m_18_), .Y(_1075_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(z_m_18_), .B(_194__bF_buf0), .Y(_1076_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1070_), .Y(_1077_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(z_m_17_), .Y(_1078_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf1), .B(_892_), .C(_1078_), .D(_244_), .Y(_1079_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(z_m_19_), .B(_234__bF_buf4), .C(_1079_), .Y(_1080_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1080_), .C(_1075_), .Y(_22__18_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1067_), .Y(_1081_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(z_m_18_), .Y(_1082_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_1082_), .Y(_1083_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(z_m_19_), .Y(_1084_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(z_m_19_), .Y(_1085_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_547_), .C(_194__bF_buf0), .D(_1085_), .Y(_1086_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(z_m_19_), .B(_1083_), .C(_1086_), .Y(_1087_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(z_m_18_), .B(_243__bF_buf0), .Y(_1088_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf1), .B(_893_), .C(_1084_), .D(_1027_), .Y(_1089_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf0), .B(z_m_20_), .C(_1089_), .Y(_1090_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_1090_), .C(_1087_), .Y(_22__19_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf1), .B(_1085_), .Y(_1091_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_1091_), .C(z_m_20_), .Y(_1092_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(z_m_20_), .Y(_1093_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf1), .B(_1093_), .C(_1085_), .Y(_1094_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(z_m_21_), .Y(_1095_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf2), .B(_894_), .C(_1095_), .D(_235_), .Y(_1096_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(z_m_19_), .B(_243__bF_buf1), .C(_1096_), .Y(_1097_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1097_), .C(_1092_), .Y(_22__20_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .Y(_1098_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(z_m_11_), .B(z_m_19_), .C(z_m_20_), .Y(_1099_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1098_), .Y(_1100_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_1100_), .C(_1082_), .Y(_1101_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1101_), .C(_1095_), .Y(_1102_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .Y(_1103_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_999_), .C(_1101_), .Y(_1104_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1105_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf4), .B(_1105_), .C(z_m_21_), .D(_548_), .Y(_1106_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(z_m_22_), .Y(_1107_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf2), .B(_895_), .C(_1107_), .D(_235_), .Y(_1108_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(z_m_20_), .B(_243__bF_buf0), .C(_1108_), .Y(_1109_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1106_), .C(_1109_), .Y(_22__21_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(z_m_22_), .B(_1104_), .Y(_1110_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .Y(_1111_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_547_), .C(_194__bF_buf0), .D(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(z_m_22_), .B(_1104_), .C(_1112_), .Y(_1113_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(z_m_21_), .B(_243__bF_buf0), .Y(_1114_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_239__bF_buf2), .B(_896_), .C(_1107_), .D(_1027_), .Y(_1115_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf4), .B(z_m_23_), .C(_1115_), .Y(_1116_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1116_), .C(_1113_), .Y(_22__22_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(z_m_19_), .B(_1082_), .Y(_1117_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1093_), .Y(_1118_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1118_), .Y(_1119_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(z_m_22_), .B(z_m_21_), .C(_1119_), .Y(_1120_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_1120_), .Y(_1121_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .B(_1121_), .Y(_1122_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .Y(_1123_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .B(_1111_), .C(state_3_bF_buf0), .Y(_1124_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .Y(_1125_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_218_), .C(_1125_), .Y(_1126_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_26_), .C(state_5_), .D(_1126_), .Y(_1127_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_224_), .C(z_m_23_), .Y(_1128_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1127_), .Y(_1129_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1124_), .B(_1123_), .C(_1129_), .Y(_22__23_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_114_), .C(_529_), .Y(_1130_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_250_), .Y(_1131_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_536_), .C(_120_), .Y(_1132_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_1131_), .C(_1132_), .Y(_1133_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1133_), .C(state_12_bF_buf0), .Y(_1134_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(z_23_), .B(_38__bF_buf1), .Y(_1135_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_221_), .Y(_1136_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1125_), .C(z_e_0_), .Y(_1137_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1137_), .C(state_11_bF_buf2), .Y(_1138_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1138_), .C(_1134_), .Y(_20__23_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_1131_), .C(_1132_), .Y(_1139_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1139_), .C(state_12_bF_buf1), .Y(_1140_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(z_24_), .B(_38__bF_buf1), .Y(_1141_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(z_e_0_), .B(_206_), .Y(_1142_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_1142_), .Y(_1143_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1143_), .C(state_11_bF_buf2), .Y(_1144_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1144_), .C(_1140_), .Y(_20__24_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_1131_), .C(_1132_), .Y(_1145_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1145_), .C(state_12_bF_buf1), .Y(_1146_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(z_25_), .B(_38__bF_buf1), .Y(_1147_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(z_e_0_), .B(z_e_1_), .Y(_1148_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .Y(_1149_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(z_e_2_), .Y(_1150_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(z_e_0_), .B(z_e_1_), .C(z_e_2_), .Y(_1151_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1150_), .Y(_1152_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_1152_), .C(state_11_bF_buf2), .Y(_1153_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1153_), .C(_1146_), .Y(_20__25_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_1131_), .C(_1132_), .Y(_1154_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1154_), .C(state_12_bF_buf0), .Y(_1155_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(z_26_), .B(_38__bF_buf1), .Y(_1156_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(z_e_2_), .B(_1149_), .C(z_e_3_), .Y(_1157_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .B(_1150_), .Y(_1158_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .Y(_1159_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1159_), .Y(_1160_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1160_), .C(state_11_bF_buf2), .Y(_1161_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .B(_1161_), .C(_1155_), .Y(_20__26_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_1131_), .C(_1132_), .Y(_1162_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1162_), .C(state_12_bF_buf0), .Y(_1163_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(z_27_), .B(_38__bF_buf2), .Y(_1164_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_1158_), .Y(_1165_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .B(_1150_), .C(z_e_4_), .Y(_1166_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1165_), .Y(_1167_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1167_), .C(state_11_bF_buf2), .Y(_1168_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1168_), .C(_1163_), .Y(_20__27_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_1131_), .C(_1132_), .Y(_1169_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1169_), .C(state_12_bF_buf0), .Y(_1170_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(z_28_), .B(_38__bF_buf2), .Y(_1171_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(z_e_4_), .B(_1159_), .C(z_e_5_), .Y(_1172_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_1159_), .C(_1172_), .Y(_1173_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1173_), .C(state_11_bF_buf2), .Y(_1174_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1174_), .C(_1170_), .Y(_20__28_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_1131_), .C(_1132_), .Y(_1175_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1175_), .C(state_12_bF_buf0), .Y(_1176_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(z_29_), .B(_38__bF_buf2), .Y(_1177_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_210_), .Y(_1178_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(z_e_6_), .Y(_1179_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf0), .B(_1179_), .C(state_11_bF_buf2), .Y(_1180_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1180_), .C(_1176_), .Y(_20__29_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_1131_), .C(_1132_), .Y(_1181_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1181_), .C(state_12_bF_buf1), .Y(_1182_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(z_30_), .B(_38__bF_buf1), .Y(_1183_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(z_e_7_), .Y(_1184_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(z_e_6_), .B(_1178_), .Y(_1185_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1185_), .Y(_1186_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(z_e_6_), .B(_1178_), .C(z_e_7_), .Y(_1187_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1186_), .Y(_1188_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .Y(_1189_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_36__bF_buf1), .B(_1189_), .C(state_11_bF_buf0), .Y(_1190_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1182_), .C(_1190_), .Y(_20__30_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_533_), .Y(_1191_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_51_), .C(z_31_), .Y(_1192_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_1131_), .C(_1192_), .Y(_1193_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_326_), .C(_536_), .Y(_1194_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(_536_), .C(_1194_), .Y(_1195_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_1191_), .C(_122_), .D(_1195_), .Y(_1196_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_1196_), .C(state_12_bF_buf2), .Y(_1197_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(state_11_bF_buf0), .B(z_s), .C(z_31_), .D(_38__bF_buf1), .Y(_1198_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1197_), .Y(_20__31_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_123_), .C(_195_), .Y(_1199_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_1200_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_1200_), .C(_899_), .Y(_1201_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1199_), .Y(_1202_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_54_), .C(_1202_), .Y(_6__23_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(dividend_0_), .Y(_1203_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_562__bF_buf5), .Y(_9__0_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(dividend_1_), .Y(_1204_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1203_), .C(_1204_), .D(_562__bF_buf5), .Y(_9__1_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(dividend_2_), .Y(_1205_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1204_), .C(_1205_), .D(_562__bF_buf5), .Y(_9__2_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(dividend_3_), .Y(_1206_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1205_), .C(_1206_), .D(_562__bF_buf5), .Y(_9__3_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(dividend_4_), .Y(_1207_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1206_), .C(_1207_), .D(_562__bF_buf5), .Y(_9__4_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(dividend_5_), .Y(_1208_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1207_), .C(_1208_), .D(_562__bF_buf6), .Y(_9__5_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(dividend_6_), .Y(_1209_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1208_), .C(_1209_), .D(_562__bF_buf3), .Y(_9__6_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(dividend_7_), .Y(_1210_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1209_), .C(_1210_), .D(_562__bF_buf3), .Y(_9__7_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(dividend_8_), .Y(_1211_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1210_), .C(_1211_), .D(_562__bF_buf5), .Y(_9__8_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(dividend_9_), .Y(_1212_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1211_), .C(_1212_), .D(_562__bF_buf5), .Y(_9__9_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(dividend_10_), .Y(_1213_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf1), .B(_1212_), .C(_1213_), .D(_562__bF_buf5), .Y(_9__10_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(dividend_11_), .Y(_1214_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1213_), .C(_1214_), .D(_562__bF_buf3), .Y(_9__11_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(dividend_12_), .Y(_1215_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1214_), .C(_1215_), .D(_562__bF_buf3), .Y(_9__12_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(dividend_13_), .Y(_1216_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1215_), .C(_1216_), .D(_562__bF_buf3), .Y(_9__13_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(dividend_14_), .Y(_1217_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1216_), .C(_1217_), .D(_562__bF_buf3), .Y(_9__14_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(dividend_15_), .Y(_1218_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf3), .B(_1217_), .C(_1218_), .D(_562__bF_buf3), .Y(_9__15_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(dividend_16_), .Y(_1219_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1218_), .C(_1219_), .D(_562__bF_buf6), .Y(_9__16_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(dividend_17_), .Y(_1220_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1219_), .C(_1220_), .D(_562__bF_buf6), .Y(_9__17_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(dividend_18_), .Y(_1221_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1220_), .C(_1221_), .D(_562__bF_buf6), .Y(_9__18_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(dividend_19_), .Y(_1222_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1221_), .C(_1222_), .D(_562__bF_buf6), .Y(_9__19_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(dividend_20_), .Y(_1223_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1222_), .C(_1223_), .D(_562__bF_buf6), .Y(_9__20_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(dividend_21_), .Y(_1224_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf0), .B(_1223_), .C(_1224_), .D(_562__bF_buf6), .Y(_9__21_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(dividend_22_), .Y(_1225_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_1224_), .C(_1225_), .D(_562__bF_buf6), .Y(_9__22_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(dividend_23_), .Y(_1226_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_1225_), .C(_1226_), .D(_562__bF_buf1), .Y(_9__23_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(dividend_24_), .Y(_1227_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_1226_), .C(_1227_), .D(_562__bF_buf1), .Y(_9__24_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(dividend_25_), .Y(_1228_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf4), .B(_1227_), .C(_1228_), .D(_562__bF_buf1), .Y(_9__25_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(dividend_26_), .B(_561__bF_buf4), .Y(_1229_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_199__bF_buf5), .B(_1228_), .C(_1229_), .Y(_9__26_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(dividend_27_), .Y(_1230_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf5), .B(a_m_0_), .C(state_14_bF_buf7), .D(dividend_26_), .Y(_1231_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_562__bF_buf4), .C(_1231_), .Y(_9__27_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(a_m_1_), .Y(_1232_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(dividend_27_), .C(dividend_28_), .D(_561__bF_buf0), .Y(_1233_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf6), .B(_1232_), .C(_1233_), .Y(_9__28_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_28_), .C(dividend_29_), .D(_561__bF_buf0), .Y(_1234_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_182__bF_buf1), .C(_1234_), .Y(_9__29_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_29_), .C(dividend_30_), .D(_561__bF_buf0), .Y(_1235_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1968_), .B(_182__bF_buf5), .C(_1235_), .Y(_9__30_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_30_), .C(dividend_31_), .D(_561__bF_buf3), .Y(_1236_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_182__bF_buf1), .C(_1236_), .Y(_9__31_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_31_), .C(dividend_32_), .D(_561__bF_buf3), .Y(_1237_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_182__bF_buf1), .C(_1237_), .Y(_9__32_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_32_), .C(dividend_33_), .D(_561__bF_buf3), .Y(_1238_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_182__bF_buf1), .C(_1238_), .Y(_9__33_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_33_), .C(dividend_34_), .D(_561__bF_buf4), .Y(_1239_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_182__bF_buf1), .C(_1239_), .Y(_9__34_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(dividend_34_), .C(dividend_35_), .D(_561__bF_buf2), .Y(_1240_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1984_), .B(_182__bF_buf6), .C(_1240_), .Y(_9__35_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_35_), .C(dividend_36_), .D(_561__bF_buf2), .Y(_1241_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_182__bF_buf6), .C(_1241_), .Y(_9__36_) );
AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_36_), .C(dividend_37_), .D(_561__bF_buf2), .Y(_1242_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1988_), .B(_182__bF_buf6), .C(_1242_), .Y(_9__37_) );
AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_37_), .C(dividend_38_), .D(_561__bF_buf1), .Y(_1243_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_182__bF_buf0), .C(_1243_), .Y(_9__38_) );
AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_38_), .C(dividend_39_), .D(_561__bF_buf1), .Y(_1244_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_182__bF_buf0), .C(_1244_), .Y(_9__39_) );
AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_39_), .C(dividend_40_), .D(_561__bF_buf1), .Y(_1245_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(_182__bF_buf0), .C(_1245_), .Y(_9__40_) );
AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_40_), .C(dividend_41_), .D(_561__bF_buf1), .Y(_1246_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_182__bF_buf0), .C(_1246_), .Y(_9__41_) );
AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_41_), .C(dividend_42_), .D(_561__bF_buf1), .Y(_1247_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_182__bF_buf0), .C(_1247_), .Y(_9__42_) );
AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_42_), .C(dividend_43_), .D(_561__bF_buf2), .Y(_1248_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .B(_182__bF_buf0), .C(_1248_), .Y(_9__43_) );
AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf4), .B(dividend_43_), .C(dividend_44_), .D(_561__bF_buf2), .Y(_1249_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_182__bF_buf6), .C(_1249_), .Y(_9__44_) );
AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(dividend_44_), .C(dividend_45_), .D(_561__bF_buf4), .Y(_1250_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_182__bF_buf6), .C(_1250_), .Y(_9__45_) );
AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(dividend_45_), .C(dividend_46_), .D(_561__bF_buf4), .Y(_1251_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_182__bF_buf6), .C(_1251_), .Y(_9__46_) );
AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_46_), .C(dividend_47_), .D(_561__bF_buf0), .Y(_1252_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_182__bF_buf1), .C(_1252_), .Y(_9__47_) );
AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_47_), .C(dividend_48_), .D(_561__bF_buf3), .Y(_1253_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_182__bF_buf1), .C(_1253_), .Y(_9__48_) );
AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(dividend_48_), .C(dividend_49_), .D(_561__bF_buf3), .Y(_1254_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_182__bF_buf5), .C(_1254_), .Y(_9__49_) );
AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf1), .B(dividend_49_), .C(dividend_50_), .D(_561__bF_buf0), .Y(_1255_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_182__bF_buf5), .C(_1255_), .Y(_9__50_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_868_), .Y(_1256_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_870_), .Y(_1257_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_861_), .B(_1256_), .C(_1257_), .Y(_1258_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(remainder_0_), .B(_253_), .Y(_1259_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1259_), .B(_667_), .Y(_1260_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1258__bF_buf5), .B(_567__bF_buf4), .C(_1260_), .Y(_1261_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(remainder_0_), .B(_871__bF_buf5), .C(state_1_bF_buf6), .Y(_1262_) );
AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(dividend_50_), .C(remainder_0_), .D(_563__bF_buf4), .Y(_1263_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1262_), .C(_1263_), .Y(_13__0_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(_222_), .Y(_1264_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(round_bit), .Y(_1265_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(sticky), .B(_1265_), .C(state_13_), .Y(_1266_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(sticky), .C(state_9_), .Y(_1267_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(_560_), .Y(_1268_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(remainder_50_), .B(remainder_49_), .Y(_1269_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_572_), .C(_1269_), .Y(_1270_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1270_), .Y(_1271_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(remainder_42_), .B(remainder_41_), .Y(_1272_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_621_), .C(_1272_), .Y(_1273_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(remainder_46_), .B(remainder_45_), .Y(_1274_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_592_), .C(_1274_), .Y(_1275_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1273_), .Y(_1276_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(remainder_34_), .B(remainder_33_), .Y(_1277_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_755_), .C(_1277_), .Y(_1278_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(remainder_38_), .B(remainder_37_), .Y(_1279_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_644_), .C(_1279_), .Y(_1280_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1280_), .Y(_1281_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1271_), .B(_1281_), .C(_1276_), .Y(_1282_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(remainder_10_), .B(remainder_9_), .Y(_1283_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_680_), .C(_1283_), .Y(_1284_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(remainder_14_), .B(remainder_13_), .Y(_1285_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_721_), .C(_1285_), .Y(_1286_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1286_), .Y(_1287_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(remainder_0_), .B(remainder_2_), .Y(_1288_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_1288_), .Y(_1289_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(remainder_6_), .B(remainder_5_), .Y(_1290_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_671_), .C(_1290_), .Y(_1291_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1291_), .Y(_1292_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(_1292_), .Y(_1293_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(remainder_26_), .B(remainder_25_), .Y(_1294_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_779_), .C(_1294_), .Y(_1295_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(remainder_30_), .B(remainder_29_), .Y(_1296_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_831_), .C(_1296_), .Y(_1297_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1297_), .Y(_1298_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(remainder_18_), .B(remainder_17_), .Y(_1299_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_705_), .C(_1299_), .Y(_1300_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(remainder_22_), .B(remainder_21_), .Y(_1301_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_791_), .C(_1301_), .Y(_1302_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1302_), .Y(_1303_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1303_), .C(_1293_), .Y(_1304_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1304_), .Y(_1305_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1305_), .C(_1266_), .Y(_19_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf0), .B(guard), .C(round_bit), .Y(_1306_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(state_13_), .B(guard), .C(_546_), .Y(_1307_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(_545_), .Y(_1308_) );
AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_1_), .C(round_bit), .D(_1308_), .Y(_1309_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1307_), .C(_1309_), .Y(_14_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_546_), .C(guard), .Y(_1310_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(z_m_0_), .B(_234__bF_buf1), .Y(_1311_) );
AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(state_9_), .B(quotient_2_), .C(round_bit), .D(_243__bF_buf2), .Y(_1312_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .B(_1311_), .C(_1312_), .Y(_11_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(a_e_0_), .B(_116_), .Y(_1313_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(a_e_0_), .Y(_1314_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(b_e_0_), .B(_1314_), .Y(_1315_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1315_), .C(state_6_bF_buf3), .Y(_1316_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(z_m_23_), .B(z_m_22_), .C(_1104_), .Y(_1317_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .Y(_1318_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf3), .B(state_3_bF_buf1), .Y(_1319_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_1319_), .Y(_1320_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .Y(_1321_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_546_), .Y(_1322_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf2), .B(_1318_), .C(_1322_), .Y(_1323_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_222_), .C(_205_), .Y(_1324_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_243__bF_buf0), .Y(_1325_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf2), .B(_1317_), .C(_1325_), .Y(_1326_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_1323_), .C(_1326_), .Y(_1327_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1327_), .Y(_21__0_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1328_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(_1122_), .Y(_1329_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(z_e_1_), .B(_1123_), .C(state_3_bF_buf3), .Y(_1330_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_546_), .C(z_e_1_), .Y(_1331_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .Y(_1332_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(_115_), .Y(_1333_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(_87_), .Y(_1334_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1334_), .Y(_1335_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1332_), .Y(_1336_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1335_), .C(state_6_bF_buf3), .Y(_1337_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1337_), .C(_1328_), .D(_244_), .Y(_1338_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf3), .B(_1328_), .C(_1338_), .Y(_1339_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1331_), .Y(_1340_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1330_), .C(_1340_), .Y(_21__1_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(z_e_2_), .B(_207_), .Y(_1341_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .Y(_1342_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(z_e_2_), .B(_207_), .Y(_1343_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1342_), .Y(_1344_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_1122_), .Y(_1345_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(z_e_2_), .B(_1123_), .C(state_3_bF_buf3), .Y(_1346_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .Y(_1347_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_234__bF_buf3), .Y(_1348_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(_1336_), .Y(_1349_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(a_e_2_), .B(b_e_2_), .Y(_1350_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .Y(_1351_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_1351_), .C(_182__bF_buf4), .Y(_1352_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_1351_), .C(_1352_), .Y(_1353_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_243__bF_buf3), .Y(_1354_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1353_), .C(_1354_), .Y(_1355_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(z_e_2_), .C(_1355_), .Y(_1356_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1346_), .C(_1356_), .Y(_21__2_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .Y(_1357_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1341_), .Y(_1358_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .B(_1342_), .Y(_1359_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1359_), .Y(_1360_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1122_), .Y(_1361_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(z_e_3_), .B(_1123_), .C(state_3_bF_buf3), .Y(_1362_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_234__bF_buf3), .Y(_1363_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(b_e_2_), .Y(_1364_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(a_e_2_), .B(_1364_), .Y(_1365_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(_1349_), .C(_1365_), .Y(_1366_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .Y(_1367_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(b_e_3_), .Y(_1368_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(a_e_3_), .B(_1368_), .Y(_1369_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(a_e_3_), .Y(_1370_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(b_e_3_), .B(_1370_), .Y(_1371_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1371_), .C(_1367_), .Y(_1372_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .Y(_1373_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .Y(_1374_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1374_), .C(_1366_), .Y(_1375_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf3), .B(_1375_), .C(_1372_), .Y(_1376_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_243__bF_buf3), .Y(_1377_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1376_), .C(_1377_), .Y(_1378_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(z_e_3_), .C(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_1362_), .C(_1379_), .Y(_21__3_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(z_e_4_), .B(_1123_), .Y(_1380_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(z_e_4_), .B(_1358_), .Y(_1381_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1341_), .C(_209_), .Y(_1382_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1381_), .Y(_1383_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_1383_), .Y(_1384_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1122_), .C(state_3_bF_buf3), .Y(_1385_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(a_e_4_), .Y(_1386_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(b_e_4_), .B(_1386_), .Y(_1387_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(b_e_4_), .B(_1386_), .Y(_1388_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .Y(_1389_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_1387_), .Y(_1390_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .Y(_1391_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1373_), .C(_1371_), .Y(_1392_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(_1391_), .Y(_1393_) );
AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_234__bF_buf3), .B(_1384_), .C(_1167_), .D(_243__bF_buf3), .Y(_1394_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf4), .B(_1393_), .C(_1394_), .Y(_1395_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(z_e_4_), .B(_1347_), .C(_1395_), .Y(_1396_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1380_), .C(_1396_), .Y(_21__4_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_1381_), .Y(_1397_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_1317_), .C(_208_), .Y(_1398_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf3), .B(_1398_), .Y(_1399_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .Y(_1400_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(z_e_5_), .B(_1400_), .C(_234__bF_buf3), .Y(_1401_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1401_), .C(_1397_), .Y(_1402_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1392_), .C(_1389_), .Y(_1403_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(a_e_5_), .Y(_1404_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(b_e_5_), .B(_1404_), .Y(_1405_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(b_e_5_), .B(_1404_), .Y(_1406_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .Y(_1407_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1405_), .Y(_1408_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1408_), .Y(_1409_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1403_), .C(state_6_bF_buf3), .Y(_1410_) );
AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf3), .B(_1173_), .C(z_e_5_), .D(_1323_), .Y(_1411_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1410_), .C(_1411_), .Y(_1412_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1402_), .Y(_21__5_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1409_), .Y(_1413_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(a_e_6_), .B(_41_), .Y(_1414_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(b_e_6_), .B(_83_), .Y(_1415_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1415_), .Y(_1416_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .Y(_1417_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(_1417_), .C(_182__bF_buf4), .Y(_1418_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(_1417_), .C(_1418_), .Y(_1419_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .Y(_1420_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1317_), .C(_211_), .Y(_1421_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .Y(_1422_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(z_e_6_), .B(_1397_), .C(_234__bF_buf3), .Y(_1423_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf2), .B(_1422_), .C(_1423_), .Y(_1424_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_1420_), .C(_1424_), .Y(_1425_) );
AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf3), .B(_1179_), .C(z_e_6_), .D(_1323_), .Y(_1426_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_1426_), .C(_1425_), .Y(_21__6_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(a_e_7_), .B(b_e_7_), .Y(_1427_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1427_), .Y(_1428_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1413_), .C(_1428_), .Y(_1429_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1413_), .Y(_1430_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1430_), .C(_1427_), .Y(_1431_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(state_6_bF_buf3), .B(_1429_), .C(_1431_), .Y(_1432_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1318_), .Y(_1433_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(z_e_6_), .B(z_e_7_), .C(_1397_), .Y(_1434_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_1420_), .C(_1184_), .Y(_1435_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1435_), .Y(_1436_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1317_), .Y(_1437_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1437_), .B(_1433_), .C(state_3_bF_buf0), .Y(_1438_) );
OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_1436_), .C(_1189_), .D(_244_), .Y(_1439_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(z_e_7_), .C(_1439_), .Y(_1440_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1440_), .C(_1432_), .Y(_21__7_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1427_), .Y(_1441_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1408_), .C(_1441_), .Y(_1442_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(b_e_7_), .Y(_1443_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(a_e_7_), .Y(_1444_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1415_), .C(_1444_), .Y(_1445_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1446_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_1446_), .C(_1407_), .Y(_1447_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1447_), .Y(_1448_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(_1445_), .Y(_1449_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1392_), .C(_1449_), .Y(_1450_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(a_e_8_), .B(b_e_8_), .Y(_1451_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1392_), .Y(_1452_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .Y(_1453_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1452_), .C(_1451_), .Y(_1454_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .Y(_1455_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_182__bF_buf4), .B(_1455_), .Y(_1456_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1451_), .C(_1456_), .Y(_1457_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf0), .B(_234__bF_buf4), .C(z_e_8_), .Y(_1458_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(state_3_bF_buf0), .C(_234__bF_buf4), .Y(_1459_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1459_), .C(_1458_), .Y(_1460_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_1434_), .C(_1460_), .Y(_1461_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_242_), .C(z_e_8_), .Y(_1462_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_242_), .Y(_1463_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_1463_), .Y(_1464_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1464_), .Y(_1465_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_224_), .Y(_1466_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_194__bF_buf2), .B(_1318_), .C(_1466_), .Y(_1467_) );
AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_1465_), .C(z_e_8_), .D(_1467_), .Y(_1468_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .B(_1468_), .C(_1461_), .Y(_21__8_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(b_e_8_), .C(_1454_), .Y(_1469_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(a_e_9_), .B(b_e_9_), .Y(_1470_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .C(_182__bF_buf4), .Y(_1471_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .C(_1471_), .Y(_1472_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_1434_), .Y(_1473_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(z_e_9_), .B(_1473_), .C(_1318_), .Y(_1474_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .Y(_1475_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1475_), .B(_1317_), .C(_34_), .Y(_1476_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(state_3_bF_buf0), .B(_1476_), .C(_1474_), .Y(_1477_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_1320_), .Y(_1478_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_1464_), .Y(_1479_) );
AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(z_e_9_), .B(_1478_), .C(state_5_), .D(_1479_), .Y(_1480_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1472_), .C(_1477_), .Y(_21__9_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_79_), .C(_531_), .Y(_1481_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_535_), .Y(_1482_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf3), .B(b_e_0_), .Y(_1483_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(b_e_0_), .B(_238_), .Y(_1484_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1485_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(b_23_), .C(_1485_), .Y(_1486_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf3), .B(_1200_), .C(_198_), .Y(_1487_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(b_e_0_), .C(_1486_), .Y(_1488_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1482_), .C(_1488_), .Y(_5__0_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(_1482_), .C(state_12_bF_buf3), .Y(_1489_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(b_m_23_), .B(b_e_0_), .Y(_1490_) );
OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_1490_), .C(state_12_bF_buf3), .D(_1200_), .Y(_1491_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_380_), .Y(_1492_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_1492_), .Y(_1493_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(b_23_), .B(b_24_), .C(_1493_), .Y(_1494_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(_1485_), .C(_1494_), .Y(_1495_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(_1491_), .C(_1495_), .Y(_1496_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1489_), .Y(_5__1_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(b_e_0_), .C(state_10_), .Y(_1497_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .Y(_1498_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf6), .B(state_10_), .C(_899_), .Y(_1499_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .Y(_1500_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .C(_1500_), .Y(_1501_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1498_), .B(_1501_), .C(b_e_2_), .Y(_1502_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(b_25_), .C(_193_), .Y(_1503_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(b_25_), .B(_1492_), .C(_1503_), .Y(_1504_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(b_e_1_), .B(b_e_2_), .Y(_1505_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1484_), .Y(_1506_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_1506_), .C(_1502_), .Y(_5__2_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(b_25_), .B(_1492_), .Y(_1507_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_1507_), .Y(_1508_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_1507_), .Y(_1509_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1510_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf3), .B(_1508_), .C(_1510_), .Y(_1511_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_118_), .Y(_1512_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .Y(_1513_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1505_), .C(_1368_), .Y(_1514_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1513_), .C(state_10_), .Y(_1515_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1511_), .Y(_1516_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(_1500_), .C(_1516_), .Y(_5__3_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_1510_), .Y(_1517_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(b_27_), .B(_1509_), .C(state_4_bF_buf3), .Y(_1518_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_1513_), .C(_1500_), .Y(_1519_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(b_e_4_), .B(_1512_), .Y(_1520_) );
AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(state_10_), .B(_1520_), .C(b_e_4_), .D(_1519_), .Y(_1521_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .B(_1518_), .C(_1521_), .Y(_5__4_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .B(b_28_), .C(_193_), .Y(_1522_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(b_28_), .B(_1517_), .C(_1522_), .Y(_1523_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(b_e_4_), .B(_1512_), .C(b_e_5_), .Y(_1524_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_1512_), .C(_1524_), .Y(_1525_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(state_10_), .B(_1525_), .Y(_1526_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf4), .B(_902_), .C(b_e_5_), .Y(_1527_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1527_), .C(_1523_), .Y(_5__5_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(b_28_), .B(_1517_), .Y(_1528_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_1528_), .C(state_4_bF_buf6), .Y(_1529_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_1528_), .C(_1529_), .Y(_1530_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_39_), .Y(_1531_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1512_), .Y(_1532_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_1512_), .C(b_e_6_), .Y(_1533_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .Y(_1534_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1534_), .C(state_10_), .Y(_1535_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_1500_), .C(_1535_), .Y(_1536_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1536_), .Y(_5__6_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_1528_), .Y(_1537_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(b_30_), .B(_1537_), .Y(_1538_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(b_30_), .Y(_1539_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1539_), .C(state_4_bF_buf6), .Y(_1540_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1512_), .C(b_e_7_), .Y(_1541_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .Y(_1542_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1532_), .Y(_1543_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .Y(_1544_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1544_), .C(state_10_), .Y(_1545_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf4), .B(_902_), .C(b_e_7_), .Y(_1546_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1546_), .C(_1540_), .Y(_5__7_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_1544_), .C(_1500_), .Y(_1547_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(b_e_8_), .B(_1543_), .Y(_1548_) );
AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(state_10_), .B(_1548_), .C(b_e_8_), .D(_1547_), .Y(_1549_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(b_30_), .B(_1529_), .C(_1549_), .Y(_5__8_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(b_e_9_), .Y(_1550_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(b_e_9_), .B(_1548_), .C(state_10_), .Y(_1551_) );
AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(b_e_9_), .B(_1499_), .C(state_4_bF_buf6), .D(_1538_), .Y(_1552_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1551_), .C(_1552_), .Y(_5__9_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_250_), .Y(_1553_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_532_), .Y(_1554_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1554_), .Y(_1555_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_536_), .Y(_1556_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1556_), .B(_1555_), .C(state_12_bF_buf2), .Y(_1557_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_1969_), .Y(_1558_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .Y(_1559_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_1559_), .C(a_e_0_), .Y(_1560_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(a_e_0_), .B(_248_), .Y(_1561_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(_441_), .C(_1561_), .Y(_1562_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .B(_1562_), .C(_1557_), .Y(_1__0_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(_1554_), .Y(_1563_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_536_), .C(state_12_bF_buf2), .Y(_1564_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(a_m_23_), .B(a_e_0_), .Y(_1565_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1565_), .C(_1558_), .Y(_1566_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1567_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .Y(_1568_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_1568_), .Y(_1569_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(a_23_), .B(a_24_), .C(_1569_), .Y(_1570_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(_1567_), .C(_1570_), .Y(_1571_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(_1566_), .C(_1571_), .Y(_1572_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1563_), .C(_1572_), .Y(_1__1_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_112_), .C(_236_), .Y(_1573_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_1573_), .C(a_e_2_), .Y(_1574_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(a_25_), .C(_193_), .Y(_1575_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(a_25_), .B(_1568_), .C(_1575_), .Y(_1576_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(a_e_1_), .B(a_e_2_), .Y(_1577_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1561_), .Y(_1578_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .B(_1578_), .C(_1574_), .Y(_1__2_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_1579_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(a_25_), .B(_1568_), .Y(_1580_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_1580_), .Y(_1581_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_1580_), .Y(_1582_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1583_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf6), .B(_1581_), .C(_1583_), .Y(_1584_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_113_), .Y(_1585_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .Y(_1586_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1577_), .C(_1370_), .Y(_1587_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(_1586_), .C(state_2_), .Y(_1588_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_1584_), .B(_1588_), .Y(_1589_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1579_), .C(_1589_), .Y(_1__3_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_1583_), .Y(_1590_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_1590_), .Y(_1591_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(a_27_), .B(_1582_), .C(_1591_), .Y(_1592_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1586_), .Y(_1593_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(a_e_4_), .B(_1585_), .Y(_1594_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(_1593_), .C(state_2_), .Y(_1595_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf4), .B(_1969_), .C(a_e_4_), .Y(_1596_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .B(_1596_), .C(_1592_), .Y(_1__4_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(a_28_), .B(_1590_), .Y(_1597_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .Y(_1598_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_1598_), .Y(_1599_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(a_28_), .B(_1590_), .C(_1599_), .Y(_1600_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1594_), .C(_1579_), .Y(_1601_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(a_e_5_), .B(_1601_), .Y(_1602_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_1585_), .Y(_1603_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_1603_), .Y(_1604_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1604_), .C(_1600_), .Y(_1__5_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_1597_), .Y(_1605_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_1605_), .Y(_1606_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(a_29_), .B(_1598_), .C(_1606_), .Y(_1607_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_81_), .Y(_1608_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1585_), .Y(_1609_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .Y(_1610_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_1603_), .C(_1610_), .Y(_1611_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_1611_), .Y(_1612_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf4), .B(_1969_), .C(a_e_6_), .Y(_1613_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1613_), .C(_1607_), .Y(_1__6_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(a_30_), .B(_1605_), .Y(_1614_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .B(a_30_), .Y(_1615_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1615_), .C(state_4_bF_buf6), .Y(_1616_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1585_), .C(a_e_7_), .Y(_1617_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .Y(_1618_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(a_e_7_), .B(_1610_), .Y(_1619_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1619_), .C(state_2_), .Y(_1620_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(state_12_bF_buf4), .B(_1969_), .C(a_e_7_), .Y(_1621_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_1621_), .C(_1616_), .Y(_1__7_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_1606_), .Y(_1622_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1619_), .C(_1579_), .Y(_1623_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(_111_), .Y(_1624_) );
AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1624_), .B(state_2_), .C(a_e_8_), .D(_1623_), .Y(_1625_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1622_), .Y(_1__8_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1624_), .C(_1579_), .Y(_1626_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(a_e_9_), .B(_1626_), .Y(_1627_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_110_), .C(_1624_), .Y(_1628_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .B(_1627_), .C(_1622_), .Y(_1__9_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_669_), .C(_667_), .Y(_1629_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(remainder_0_), .B(_253_), .Y(_1630_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(remainder_1_), .B(_255_), .Y(_1631_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_666_), .C(_1630_), .Y(_1632_) );
AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1632_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1633_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(remainder_1_), .B(_871__bF_buf5), .C(state_1_bF_buf4), .Y(_1634_) );
AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_0_), .C(remainder_1_), .D(_563__bF_buf6), .Y(_1635_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_1634_), .C(_1635_), .Y(_13__1_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1630_), .B(_1631_), .C(_665_), .Y(_1636_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_1636_), .Y(_1637_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_677_), .Y(_1638_) );
AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1638_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1639_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(remainder_2_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1640_) );
AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_1_), .C(remainder_2_), .D(_563__bF_buf6), .Y(_1641_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1640_), .C(_1641_), .Y(_13__2_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(divisor_2_), .B(_673_), .C(_1637_), .Y(_1642_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1642_), .B(_675_), .Y(_1643_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf1), .B(_1643_), .Y(_1644_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(remainder_3_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1645_) );
AOI22X1 AOI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_2_), .C(remainder_3_), .D(_563__bF_buf6), .Y(_1646_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_1645_), .C(_1646_), .Y(_13__3_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(divisor_4_), .B(remainder_4_), .Y(_1647_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_679_), .Y(_1648_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(_1647_), .Y(_1649_) );
AOI22X1 AOI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1649_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1650_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(remainder_4_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1651_) );
AOI22X1 AOI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_3_), .C(remainder_4_), .D(_563__bF_buf6), .Y(_1652_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1651_), .C(_1652_), .Y(_13__4_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(divisor_4_), .B(_692_), .C(_1648_), .Y(_1653_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_694_), .Y(_1654_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf1), .B(_1654_), .Y(_1655_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(remainder_5_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1656_) );
AOI22X1 AOI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_4_), .C(remainder_5_), .D(_563__bF_buf6), .Y(_1657_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1656_), .C(_1657_), .Y(_13__5_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(_695_), .Y(_1658_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(_701_), .C(_1658_), .Y(_1659_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_697_), .Y(_1660_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_1659_), .Y(_1661_) );
AOI22X1 AOI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1661_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1662_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(remainder_6_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1663_) );
AOI22X1 AOI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_5_), .C(remainder_6_), .D(_563__bF_buf6), .Y(_1664_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1662_), .B(_1663_), .C(_1664_), .Y(_13__6_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(divisor_6_), .B(_682_), .C(_1660_), .Y(_1665_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_686_), .Y(_1666_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf5), .B(_1666_), .Y(_1667_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(remainder_7_), .B(_871__bF_buf5), .C(state_1_bF_buf4), .Y(_1668_) );
AOI22X1 AOI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_6_), .C(remainder_7_), .D(_563__bF_buf6), .Y(_1669_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1668_), .C(_1669_), .Y(_13__7_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_703_), .Y(_1670_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_729_), .Y(_1671_) );
AOI22X1 AOI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1670_), .B(_1671_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1672_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(remainder_8_), .B(_871__bF_buf5), .C(state_1_bF_buf4), .Y(_1673_) );
AOI22X1 AOI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_7_), .C(remainder_8_), .D(_563__bF_buf6), .Y(_1674_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .B(_1673_), .C(_1674_), .Y(_13__8_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_726_), .Y(_1675_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .B(_730_), .Y(_1676_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf5), .B(_1676_), .Y(_1677_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(remainder_9_), .B(_871__bF_buf1), .C(state_1_bF_buf4), .Y(_1678_) );
AOI22X1 AOI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf2), .B(remainder_8_), .C(remainder_9_), .D(_563__bF_buf4), .Y(_1679_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1677_), .B(_1678_), .C(_1679_), .Y(_13__9_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_675_), .C(_1636_), .Y(_1680_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_701_), .Y(_1681_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_1680_), .C(_1681_), .Y(_1682_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_1682_), .C(_731_), .Y(_1683_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_1683_), .Y(_1684_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_1684_), .Y(_1685_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1684_), .B(_735_), .Y(_1686_) );
AOI22X1 AOI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_1686_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1687_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(remainder_10_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1688_) );
AOI22X1 AOI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_9_), .C(remainder_10_), .D(_563__bF_buf4), .Y(_1689_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1688_), .C(_1689_), .Y(_13__10_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(divisor_10_), .B(_740_), .C(_1685_), .Y(_1690_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .B(_723_), .Y(_1691_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf6), .B(_1691_), .Y(_1692_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(remainder_11_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1693_) );
AOI22X1 AOI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_10_), .C(remainder_11_), .D(_563__bF_buf4), .Y(_1694_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1693_), .C(_1694_), .Y(_13__11_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(_713_), .Y(_1695_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(_744_), .Y(_1696_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_703_), .C(_1696_), .Y(_1697_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1695_), .Y(_1698_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1697_), .Y(_1699_) );
AOI22X1 AOI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1699_), .C(_567__bF_buf4), .D(_1258__bF_buf5), .Y(_1700_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(remainder_12_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1701_) );
AOI22X1 AOI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_11_), .C(remainder_12_), .D(_563__bF_buf4), .Y(_1702_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1700_), .B(_1701_), .C(_1702_), .Y(_13__12_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(divisor_12_), .B(_711_), .C(_1699_), .Y(_1703_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_717_), .Y(_1704_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf5), .B(_1704_), .Y(_1705_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(remainder_13_), .B(_871__bF_buf5), .C(state_1_bF_buf6), .Y(_1706_) );
AOI22X1 AOI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_12_), .C(remainder_13_), .D(_563__bF_buf4), .Y(_1707_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1706_), .C(_1707_), .Y(_13__13_) );
AOI22X1 AOI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_746_), .C(_718_), .D(_1697_), .Y(_1708_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1708_), .B(_708_), .Y(_1709_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_1708_), .Y(_1710_) );
AOI22X1 AOI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(_1710_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1711_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(remainder_14_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1712_) );
AOI22X1 AOI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_13_), .C(remainder_14_), .D(_563__bF_buf4), .Y(_1713_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1712_), .C(_1713_), .Y(_13__14_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_707_), .Y(_1714_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_749_), .Y(_1715_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_1708_), .C(_1715_), .Y(_1716_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1716_), .B(_1714_), .Y(_1717_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1716_), .Y(_1718_) );
AOI22X1 AOI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(_1718_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1719_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(remainder_15_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1720_) );
AOI22X1 AOI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_14_), .C(remainder_15_), .D(_563__bF_buf4), .Y(_1721_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_1720_), .C(_1721_), .Y(_13__15_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_719_), .Y(_1722_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_1682_), .C(_1722_), .Y(_1723_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(_752_), .C(_806_), .Y(_1724_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .Y(_1725_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_806_), .C(_1723_), .Y(_1726_) );
AOI22X1 AOI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_1726_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1727_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(remainder_16_), .B(_871__bF_buf2), .C(state_1_bF_buf3), .Y(_1728_) );
AOI22X1 AOI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_15_), .C(remainder_16_), .D(_563__bF_buf3), .Y(_1729_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1728_), .C(_1729_), .Y(_13__16_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(divisor_16_), .B(_804_), .C(_1725_), .Y(_1730_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_802_), .Y(_1731_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf2), .B(_1731_), .Y(_1732_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(remainder_17_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1733_) );
AOI22X1 AOI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_16_), .C(remainder_17_), .D(_563__bF_buf3), .Y(_1734_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1732_), .B(_1733_), .C(_1734_), .Y(_13__17_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_1724_), .C(_801_), .Y(_1735_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_797_), .Y(_1736_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_1735_), .Y(_1737_) );
AOI22X1 AOI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1737_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1738_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(remainder_18_), .B(_871__bF_buf6), .C(state_1_bF_buf6), .Y(_1739_) );
AOI22X1 AOI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf6), .B(remainder_17_), .C(remainder_18_), .D(_563__bF_buf3), .Y(_1740_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1738_), .B(_1739_), .C(_1740_), .Y(_13__18_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_1735_), .C(_794_), .Y(_1741_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(_811_), .Y(_1742_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf2), .B(_1742_), .Y(_1743_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(remainder_19_), .B(_871__bF_buf2), .C(state_1_bF_buf3), .Y(_1744_) );
AOI22X1 AOI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_18_), .C(remainder_19_), .D(_563__bF_buf3), .Y(_1745_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(_1744_), .C(_1745_), .Y(_13__19_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_808_), .C(_818_), .Y(_1746_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_1746_), .Y(_1747_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .B(_787_), .Y(_1748_) );
AOI22X1 AOI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_1748_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1749_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(remainder_20_), .B(_871__bF_buf0), .C(state_1_bF_buf3), .Y(_1750_) );
AOI22X1 AOI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_19_), .C(remainder_20_), .D(_563__bF_buf2), .Y(_1751_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(_1750_), .C(_1751_), .Y(_13__20_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_1746_), .C(_784_), .Y(_1752_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_783_), .Y(_1753_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf0), .B(_1753_), .Y(_1754_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(remainder_21_), .B(_871__bF_buf0), .C(state_1_bF_buf1), .Y(_1755_) );
AOI22X1 AOI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(remainder_20_), .C(remainder_21_), .D(_563__bF_buf2), .Y(_1756_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .B(_1755_), .C(_1756_), .Y(_13__21_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_1746_), .C(_821_), .Y(_1757_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_1757_), .Y(_1758_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(_781_), .Y(_1759_) );
AOI22X1 AOI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1759_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1760_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(remainder_22_), .B(_871__bF_buf0), .C(state_1_bF_buf1), .Y(_1761_) );
AOI22X1 AOI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(remainder_21_), .C(remainder_22_), .D(_563__bF_buf2), .Y(_1762_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1760_), .B(_1761_), .C(_1762_), .Y(_13__22_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_780_), .Y(_1763_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(divisor_22_), .B(_822_), .C(_1758_), .Y(_1764_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_1763_), .Y(_1765_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf7), .B(_1765_), .Y(_1766_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(remainder_23_), .B(_871__bF_buf7), .C(state_1_bF_buf1), .Y(_1767_) );
AOI22X1 AOI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf7), .B(remainder_22_), .C(remainder_23_), .D(_563__bF_buf2), .Y(_1768_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1766_), .B(_1767_), .C(_1768_), .Y(_13__23_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_827_), .Y(_1769_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(_752_), .C(_809_), .Y(_1770_) );
NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(_1770_), .Y(_1771_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_771_), .Y(_1772_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_1771_), .Y(_1773_) );
AOI22X1 AOI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1772_), .B(_1773_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1774_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(remainder_24_), .B(_871__bF_buf7), .C(state_1_bF_buf3), .Y(_1775_) );
AOI22X1 AOI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_23_), .C(remainder_24_), .D(_563__bF_buf2), .Y(_1776_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1775_), .C(_1776_), .Y(_13__24_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_1771_), .C(_768_), .Y(_1777_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_767_), .Y(_1778_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf0), .B(_1778_), .Y(_1779_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(remainder_25_), .B(_871__bF_buf0), .C(state_1_bF_buf3), .Y(_1780_) );
AOI22X1 AOI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_24_), .C(remainder_25_), .D(_563__bF_buf1), .Y(_1781_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .B(_1780_), .C(_1781_), .Y(_13__25_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_1771_), .C(_830_), .Y(_1782_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_1782_), .Y(_1783_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1782_), .B(_774_), .Y(_1784_) );
AOI22X1 AOI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1784_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1785_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(remainder_26_), .B(_871__bF_buf0), .C(state_1_bF_buf3), .Y(_1786_) );
AOI22X1 AOI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_25_), .C(remainder_26_), .D(_563__bF_buf2), .Y(_1787_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_1786_), .C(_1787_), .Y(_13__26_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(divisor_26_), .B(_832_), .C(_1783_), .Y(_1788_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_773_), .Y(_1789_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_1788_), .Y(_1790_) );
AOI22X1 AOI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1790_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1791_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(remainder_27_), .B(_871__bF_buf2), .C(state_1_bF_buf3), .Y(_1792_) );
AOI22X1 AOI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_26_), .C(remainder_27_), .D(_563__bF_buf1), .Y(_1793_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1791_), .B(_1792_), .C(_1793_), .Y(_13__27_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_764_), .Y(_1794_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_1795_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(_1770_), .C(_776_), .Y(_1796_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(_1796_), .Y(_1797_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_1794_), .Y(_1798_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_1797_), .Y(_1799_) );
AOI22X1 AOI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1799_), .C(_567__bF_buf5), .D(_1258__bF_buf2), .Y(_1800_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(remainder_28_), .B(_871__bF_buf2), .C(state_1_bF_buf3), .Y(_1801_) );
AOI22X1 AOI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_27_), .C(remainder_28_), .D(_563__bF_buf3), .Y(_1802_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1801_), .C(_1802_), .Y(_13__28_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_761_), .Y(_1803_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_760_), .Y(_1804_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_1803_), .Y(_1805_) );
AOI22X1 AOI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_1805_), .C(_567__bF_buf5), .D(_1258__bF_buf3), .Y(_1806_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(remainder_29_), .B(_871__bF_buf2), .C(state_1_bF_buf3), .Y(_1807_) );
AOI22X1 AOI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_28_), .C(remainder_29_), .D(_563__bF_buf3), .Y(_1808_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1806_), .B(_1807_), .C(_1808_), .Y(_13__29_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_765_), .C(_840_), .Y(_1809_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_758_), .Y(_1810_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_1809_), .Y(_1811_) );
AOI22X1 AOI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1811_), .C(_567__bF_buf1), .D(_1258__bF_buf3), .Y(_1812_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(remainder_30_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1813_) );
AOI22X1 AOI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf0), .B(remainder_29_), .C(remainder_30_), .D(_563__bF_buf3), .Y(_1814_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_1812_), .B(_1813_), .C(_1814_), .Y(_13__30_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(_836_), .Y(_1815_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_1809_), .C(_1815_), .Y(_1816_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_756_), .C(_1816_), .Y(_1817_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_1815_), .C(_1810_), .Y(_1818_) );
AOI22X1 AOI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1817_), .C(_567__bF_buf1), .D(_1258__bF_buf3), .Y(_1819_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(remainder_31_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1820_) );
AOI22X1 AOI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_30_), .C(remainder_31_), .D(_563__bF_buf5), .Y(_1821_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(_1820_), .C(_1821_), .Y(_13__31_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_845_), .Y(_1822_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_848_), .Y(_1823_) );
AOI22X1 AOI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1822_), .B(_1823_), .C(_567__bF_buf0), .D(_1258__bF_buf1), .Y(_1824_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(remainder_32_), .B(_871__bF_buf2), .C(state_1_bF_buf5), .Y(_1825_) );
AOI22X1 AOI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_31_), .C(remainder_32_), .D(_563__bF_buf5), .Y(_1826_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_1824_), .B(_1825_), .C(_1826_), .Y(_13__32_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_845_), .C(_651_), .Y(_1827_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_654_), .Y(_1828_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf7), .B(_1828_), .Y(_1829_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(remainder_33_), .B(_871__bF_buf7), .C(state_1_bF_buf1), .Y(_1830_) );
AOI22X1 AOI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_32_), .C(remainder_33_), .D(_563__bF_buf1), .Y(_1831_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(_1830_), .C(_1831_), .Y(_13__33_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(divisor_33_), .B(_652_), .C(_651_), .Y(_1832_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .Y(_1833_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_845_), .C(_1833_), .Y(_1834_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(_653_), .Y(_1835_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .Y(_1836_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_643_), .Y(_1837_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_1836_), .Y(_1838_) );
AOI22X1 AOI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1838_), .C(_567__bF_buf2), .D(_1258__bF_buf4), .Y(_1839_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(remainder_34_), .B(_871__bF_buf7), .C(state_1_bF_buf1), .Y(_1840_) );
AOI22X1 AOI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_33_), .C(remainder_34_), .D(_563__bF_buf0), .Y(_1841_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1840_), .C(_1841_), .Y(_13__34_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(_641_), .C(_656_), .Y(_1842_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_648_), .Y(_1843_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_646_), .C(_1842_), .Y(_1844_) );
AOI22X1 AOI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_1843_), .C(_567__bF_buf2), .D(_1258__bF_buf4), .Y(_1845_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(remainder_35_), .B(_871__bF_buf7), .C(state_1_bF_buf1), .Y(_1846_) );
AOI22X1 AOI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_34_), .C(remainder_35_), .D(_563__bF_buf0), .Y(_1847_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_1845_), .B(_1846_), .C(_1847_), .Y(_13__35_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(_638_), .Y(_1848_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_845_), .C(_659_), .Y(_1849_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_1848_), .Y(_1850_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1849_), .Y(_1851_) );
AOI22X1 AOI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1851_), .C(_567__bF_buf3), .D(_1258__bF_buf4), .Y(_1852_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(remainder_36_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1853_) );
AOI22X1 AOI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_35_), .C(remainder_36_), .D(_563__bF_buf0), .Y(_1854_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1853_), .C(_1854_), .Y(_13__36_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_628_), .Y(_1855_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_635_), .Y(_1856_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_1855_), .Y(_1857_) );
AOI22X1 AOI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1856_), .B(_1857_), .C(_567__bF_buf3), .D(_1258__bF_buf0), .Y(_1858_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(remainder_37_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1859_) );
AOI22X1 AOI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_36_), .C(remainder_37_), .D(_563__bF_buf0), .Y(_1860_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_1858_), .B(_1859_), .C(_1860_), .Y(_13__37_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_639_), .Y(_1861_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_1861_), .C(_632_), .Y(_1862_) );
NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_1861_), .Y(_1863_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_1863_), .Y(_1864_) );
AOI22X1 AOI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1864_), .C(_567__bF_buf2), .D(_1258__bF_buf4), .Y(_1865_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(remainder_38_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1866_) );
AOI22X1 AOI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_37_), .C(remainder_38_), .D(_563__bF_buf1), .Y(_1867_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(_1866_), .C(_1867_), .Y(_13__38_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_1863_), .C(_660_), .Y(_1868_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_1868_), .Y(_1869_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_625_), .C(_1862_), .Y(_1870_) );
AOI22X1 AOI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_567__bF_buf3), .B(_1258__bF_buf0), .C(_1870_), .D(_1869_), .Y(_1871_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(remainder_39_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1872_) );
AOI22X1 AOI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_38_), .C(remainder_39_), .D(_563__bF_buf1), .Y(_1873_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_1871_), .C(_1873_), .Y(_13__39_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_853_), .Y(_1874_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_614_), .Y(_1875_) );
AOI22X1 AOI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1874_), .B(_1875_), .C(_567__bF_buf3), .D(_1258__bF_buf0), .Y(_1876_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(remainder_40_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1877_) );
AOI22X1 AOI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_39_), .C(remainder_40_), .D(_563__bF_buf1), .Y(_1878_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_1877_), .C(_1878_), .Y(_13__40_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(divisor_40_), .B(_612_), .C(_1874_), .Y(_1879_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_610_), .Y(_1880_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_871__bF_buf4), .B(_1880_), .Y(_1881_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(remainder_41_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1882_) );
AOI22X1 AOI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_40_), .C(remainder_41_), .D(_563__bF_buf1), .Y(_1883_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(_1882_), .C(_1883_), .Y(_13__41_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_591_), .Y(_1884_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_616_), .C(_602_), .Y(_1885_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_1884_), .Y(_1886_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1884_), .B(_1885_), .Y(_1887_) );
AOI22X1 AOI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(_1887_), .C(_567__bF_buf3), .D(_1258__bF_buf0), .Y(_1888_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(remainder_42_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1889_) );
AOI22X1 AOI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_41_), .C(remainder_42_), .D(_563__bF_buf5), .Y(_1890_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(_1889_), .C(_1890_), .Y(_13__42_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_1884_), .B(_1885_), .C(_591_), .Y(_1891_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_1891_), .Y(_1892_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_595_), .Y(_1893_) );
AOI22X1 AOI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_1893_), .C(_567__bF_buf3), .D(_1258__bF_buf0), .Y(_1894_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(remainder_43_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1895_) );
AOI22X1 AOI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_42_), .C(remainder_43_), .D(_563__bF_buf5), .Y(_1896_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1895_), .C(_1896_), .Y(_13__43_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_618_), .C(_605_), .Y(_1897_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_1897_), .Y(_1898_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(_618_), .Y(_1899_) );
NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_787_), .Y(_1900_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_781_), .C(_1900_), .Y(_1901_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_807_), .Y(_1902_) );
NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1901_), .Y(_1903_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_776_), .C(_1903_), .Y(_1904_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(_752_), .C(_1904_), .Y(_1905_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_1905_), .C(_851_), .Y(_1906_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(_664_), .C(_1899_), .Y(_1907_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_1907_), .C(_585_), .Y(_1908_) );
AOI22X1 AOI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1898_), .B(_1908_), .C(_567__bF_buf1), .D(_1258__bF_buf3), .Y(_1909_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(remainder_44_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1910_) );
AOI22X1 AOI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_43_), .C(remainder_44_), .D(_563__bF_buf5), .Y(_1911_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_1909_), .B(_1910_), .C(_1911_), .Y(_13__44_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_1897_), .C(_582_), .Y(_1912_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_1912_), .Y(_1913_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_579_), .Y(_1914_) );
AOI22X1 AOI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1913_), .B(_1914_), .C(_567__bF_buf1), .D(_1258__bF_buf3), .Y(_1915_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(remainder_45_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1916_) );
AOI22X1 AOI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_44_), .C(remainder_45_), .D(_563__bF_buf5), .Y(_1917_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_1916_), .C(_1917_), .Y(_13__45_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_1897_), .C(_606_), .Y(_1918_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_1918_), .Y(_1919_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(_571_), .Y(_1920_) );
AOI22X1 AOI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1919_), .B(_1920_), .C(_567__bF_buf1), .D(_1258__bF_buf3), .Y(_1921_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(remainder_46_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1922_) );
AOI22X1 AOI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_45_), .C(remainder_46_), .D(_563__bF_buf5), .Y(_1923_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_1922_), .C(_1923_), .Y(_13__46_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(_571_), .Y(_1924_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(_586_), .Y(_1925_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_1907_), .C(_1925_), .Y(_1926_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_606_), .C(_1924_), .Y(_1927_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_1927_), .C(_575_), .Y(_1928_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(_575_), .Y(_1929_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_1929_), .C(_1919_), .Y(_1930_) );
AOI22X1 AOI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_567__bF_buf1), .B(_1258__bF_buf0), .C(_1930_), .D(_1928_), .Y(_1931_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(remainder_47_), .B(_871__bF_buf3), .C(state_1_bF_buf5), .Y(_1932_) );
AOI22X1 AOI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf3), .B(remainder_46_), .C(remainder_47_), .D(_563__bF_buf5), .Y(_1933_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1931_), .C(_1933_), .Y(_13__47_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_855_), .Y(_1934_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_609_), .Y(_1935_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_1935_), .Y(_1936_) );
AOI22X1 AOI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(_1936_), .C(_567__bF_buf2), .D(_1258__bF_buf4), .Y(_1937_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(remainder_48_), .B(_871__bF_buf4), .C(state_1_bF_buf0), .Y(_1938_) );
AOI22X1 AOI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_47_), .C(remainder_48_), .D(_563__bF_buf0), .Y(_1939_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1938_), .C(_1939_), .Y(_13__48_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_867_), .C(_1934_), .Y(_1940_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_1935_), .C(_860_), .Y(_1941_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_1941_), .Y(_1942_) );
AOI22X1 AOI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1258__bF_buf4), .B(_567__bF_buf2), .C(_1940_), .D(_1942_), .Y(_1943_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(remainder_49_), .B(_871__bF_buf7), .C(state_1_bF_buf0), .Y(_1944_) );
AOI22X1 AOI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_48_), .C(remainder_49_), .D(_563__bF_buf0), .Y(_1945_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(_1943_), .C(_1945_), .Y(_13__49_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_324_), .Y(_1946_) );
NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_565_), .Y(_1947_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_869_), .C(_1947_), .Y(_1948_) );
AOI22X1 AOI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(state_14_bF_buf5), .B(remainder_49_), .C(remainder_50_), .D(_563__bF_buf0), .Y(_1949_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1948_), .C(_1949_), .Y(_13__50_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1972_), .C(a_m_0_), .Y(_1950_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_395_), .C(_1950_), .Y(_2__0_) );
AOI22X1 AOI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf2), .B(a_1_), .C(a_m_0_), .D(_1974__bF_buf0), .Y(_1951_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1973__bF_buf2), .C(_1951_), .Y(_2__1_) );
AOI22X1 AOI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(state_4_bF_buf4), .B(a_2_), .C(a_m_1_), .D(_1974__bF_buf3), .Y(_1952_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_1973__bF_buf0), .C(_1952_), .Y(_2__2_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .Y(input_a_ack) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(input_b_ack) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_2006__0_), .Y(output_z[0]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_2006__1_), .Y(output_z[1]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_2006__2_), .Y(output_z[2]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_2006__3_), .Y(output_z[3]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_2006__4_), .Y(output_z[4]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_2006__5_), .Y(output_z[5]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_2006__6_), .Y(output_z[6]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_2006__7_), .Y(output_z[7]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_2006__8_), .Y(output_z[8]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_2006__9_), .Y(output_z[9]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_2006__10_), .Y(output_z[10]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_2006__11_), .Y(output_z[11]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_2006__12_), .Y(output_z[12]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_2006__13_), .Y(output_z[13]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_2006__14_), .Y(output_z[14]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_2006__15_), .Y(output_z[15]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_2006__16_), .Y(output_z[16]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_2006__17_), .Y(output_z[17]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_2006__18_), .Y(output_z[18]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_2006__19_), .Y(output_z[19]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_2006__20_), .Y(output_z[20]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_2006__21_), .Y(output_z[21]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_2006__22_), .Y(output_z[22]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_2006__23_), .Y(output_z[23]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_2006__24_), .Y(output_z[24]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_2006__25_), .Y(output_z[25]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_2006__26_), .Y(output_z[26]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_2006__27_), .Y(output_z[27]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_2006__28_), .Y(output_z[28]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_2006__29_), .Y(output_z[29]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_2006__30_), .Y(output_z[30]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_2006__31_), .Y(output_z[31]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .Y(output_z_stb) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_1960_), .Q(state_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_1956_), .Q(state_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_1966_), .Q(state_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1959_), .Q(state_3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_1958_), .Q(state_4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1964_), .Q(state_5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1955_), .Q(state_6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_1967_), .Q(state_7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_1965_), .Q(state_8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1957_), .Q(state_9_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1963_), .Q(state_10_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1954_), .Q(state_11_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1953_), .Q(state_12_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1962_), .Q(state_13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1961_), .Q(state_14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_18_), .Q(_2007_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17__0_), .Q(_2006__0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17__1_), .Q(_2006__1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17__2_), .Q(_2006__2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17__3_), .Q(_2006__3_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17__4_), .Q(_2006__4_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17__5_), .Q(_2006__5_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17__6_), .Q(_2006__6_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__7_), .Q(_2006__7_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17__8_), .Q(_2006__8_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17__9_), .Q(_2006__9_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17__10_), .Q(_2006__10_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17__11_), .Q(_2006__11_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17__12_), .Q(_2006__12_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17__13_), .Q(_2006__13_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17__14_), .Q(_2006__14_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17__15_), .Q(_2006__15_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17__16_), .Q(_2006__16_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17__17_), .Q(_2006__17_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17__18_), .Q(_2006__18_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17__19_), .Q(_2006__19_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17__20_), .Q(_2006__20_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17__21_), .Q(_2006__21_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17__22_), .Q(_2006__22_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__23_), .Q(_2006__23_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__24_), .Q(_2006__24_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__25_), .Q(_2006__25_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17__26_), .Q(_2006__26_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17__27_), .Q(_2006__27_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__28_), .Q(_2006__28_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17__29_), .Q(_2006__29_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17__30_), .Q(_2006__30_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17__31_), .Q(_2006__31_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_15_), .Q(_2004_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_16_), .Q(_2005_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_0__0_), .Q(a_0_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_0__1_), .Q(a_1_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__2_), .Q(a_2_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__3_), .Q(a_3_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__4_), .Q(a_4_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__5_), .Q(a_5_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_0__6_), .Q(a_6_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__7_), .Q(a_7_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__8_), .Q(a_8_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_0__9_), .Q(a_9_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_0__10_), .Q(a_10_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__11_), .Q(a_11_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_0__12_), .Q(a_12_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_0__13_), .Q(a_13_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_0__14_), .Q(a_14_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__15_), .Q(a_15_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__16_), .Q(a_16_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__17_), .Q(a_17_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_0__18_), .Q(a_18_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__19_), .Q(a_19_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_0__20_), .Q(a_20_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__21_), .Q(a_21_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__22_), .Q(a_22_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_0__23_), .Q(a_23_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_0__24_), .Q(a_24_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_0__25_), .Q(a_25_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_0__26_), .Q(a_26_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_0__27_), .Q(a_27_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_0__28_), .Q(a_28_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_0__29_), .Q(a_29_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_0__30_), .Q(a_30_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__31_), .Q(a_31_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4__0_), .Q(b_0_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4__1_), .Q(b_1_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__2_), .Q(b_2_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4__3_), .Q(b_3_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_4__4_), .Q(b_4_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__5_), .Q(b_5_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__6_), .Q(b_6_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__7_), .Q(b_7_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__8_), .Q(b_8_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_4__9_), .Q(b_9_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_4__10_), .Q(b_10_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__11_), .Q(b_11_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4__12_), .Q(b_12_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4__13_), .Q(b_13_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__14_), .Q(b_14_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4__15_), .Q(b_15_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__16_), .Q(b_16_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__17_), .Q(b_17_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4__18_), .Q(b_18_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4__19_), .Q(b_19_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4__20_), .Q(b_20_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__21_), .Q(b_21_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4__22_), .Q(b_22_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__23_), .Q(b_23_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_4__24_), .Q(b_24_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_4__25_), .Q(b_25_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4__26_), .Q(b_26_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_4__27_), .Q(b_27_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4__28_), .Q(b_28_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__29_), .Q(b_29_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_4__30_), .Q(b_30_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__31_), .Q(b_31_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_20__0_), .Q(z_0_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_20__1_), .Q(z_1_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_20__2_), .Q(z_2_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20__3_), .Q(z_3_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_20__4_), .Q(z_4_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_20__5_), .Q(z_5_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_20__6_), .Q(z_6_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20__7_), .Q(z_7_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_20__8_), .Q(z_8_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_20__9_), .Q(z_9_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20__10_), .Q(z_10_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_20__11_), .Q(z_11_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_20__12_), .Q(z_12_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_20__13_), .Q(z_13_) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_20__14_), .Q(z_14_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20__15_), .Q(z_15_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_20__16_), .Q(z_16_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_20__17_), .Q(z_17_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_20__18_), .Q(z_18_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_20__19_), .Q(z_19_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_20__20_), .Q(z_20_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_20__21_), .Q(z_21_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_20__22_), .Q(z_22_) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_20__23_), .Q(z_23_) );
DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_20__24_), .Q(z_24_) );
DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_20__25_), .Q(z_25_) );
DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_20__26_), .Q(z_26_) );
DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_20__27_), .Q(z_27_) );
DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_20__28_), .Q(z_28_) );
DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_20__29_), .Q(z_29_) );
DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_20__30_), .Q(z_30_) );
DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_20__31_), .Q(z_31_) );
DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_2__0_), .Q(a_m_0_) );
DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2__1_), .Q(a_m_1_) );
DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2__2_), .Q(a_m_2_) );
DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_2__3_), .Q(a_m_3_) );
DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__4_), .Q(a_m_4_) );
DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__5_), .Q(a_m_5_) );
DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__6_), .Q(a_m_6_) );
DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_2__7_), .Q(a_m_7_) );
DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__8_), .Q(a_m_8_) );
DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_2__9_), .Q(a_m_9_) );
DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2__10_), .Q(a_m_10_) );
DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2__11_), .Q(a_m_11_) );
DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__12_), .Q(a_m_12_) );
DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_2__13_), .Q(a_m_13_) );
DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_2__14_), .Q(a_m_14_) );
DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2__15_), .Q(a_m_15_) );
DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__16_), .Q(a_m_16_) );
DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__17_), .Q(a_m_17_) );
DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__18_), .Q(a_m_18_) );
DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__19_), .Q(a_m_19_) );
DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__20_), .Q(a_m_20_) );
DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__21_), .Q(a_m_21_) );
DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__22_), .Q(a_m_22_) );
DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_2__23_), .Q(a_m_23_) );
DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6__0_), .Q(b_m_0_) );
DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6__1_), .Q(b_m_1_) );
DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6__2_), .Q(b_m_2_) );
DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6__3_), .Q(b_m_3_) );
DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6__4_), .Q(b_m_4_) );
DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__5_), .Q(b_m_5_) );
DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6__6_), .Q(b_m_6_) );
DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6__7_), .Q(b_m_7_) );
DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6__8_), .Q(b_m_8_) );
DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6__9_), .Q(b_m_9_) );
DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6__10_), .Q(b_m_10_) );
DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6__11_), .Q(b_m_11_) );
DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__12_), .Q(b_m_12_) );
DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6__13_), .Q(b_m_13_) );
DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6__14_), .Q(b_m_14_) );
DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6__15_), .Q(b_m_15_) );
DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__16_), .Q(b_m_16_) );
DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__17_), .Q(b_m_17_) );
DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__18_), .Q(b_m_18_) );
DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__19_), .Q(b_m_19_) );
DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__20_), .Q(b_m_20_) );
DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6__21_), .Q(b_m_21_) );
DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6__22_), .Q(b_m_22_) );
DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6__23_), .Q(b_m_23_) );
DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_22__0_), .Q(z_m_0_) );
DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_22__1_), .Q(z_m_1_) );
DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_22__2_), .Q(z_m_2_) );
DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_22__3_), .Q(z_m_3_) );
DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_22__4_), .Q(z_m_4_) );
DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_22__5_), .Q(z_m_5_) );
DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__6_), .Q(z_m_6_) );
DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__7_), .Q(z_m_7_) );
DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_22__8_), .Q(z_m_8_) );
DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__9_), .Q(z_m_9_) );
DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__10_), .Q(z_m_10_) );
DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__11_), .Q(z_m_11_) );
DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__12_), .Q(z_m_12_) );
DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_22__13_), .Q(z_m_13_) );
DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__14_), .Q(z_m_14_) );
DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__15_), .Q(z_m_15_) );
DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__16_), .Q(z_m_16_) );
DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__17_), .Q(z_m_17_) );
DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__18_), .Q(z_m_18_) );
DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__19_), .Q(z_m_19_) );
DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__20_), .Q(z_m_20_) );
DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_22__21_), .Q(z_m_21_) );
DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_22__22_), .Q(z_m_22_) );
DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_22__23_), .Q(z_m_23_) );
DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1__0_), .Q(a_e_0_) );
DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1__1_), .Q(a_e_1_) );
DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1__2_), .Q(a_e_2_) );
DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1__3_), .Q(a_e_3_) );
DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1__4_), .Q(a_e_4_) );
DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1__5_), .Q(a_e_5_) );
DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1__6_), .Q(a_e_6_) );
DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1__7_), .Q(a_e_7_) );
DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1__8_), .Q(a_e_8_) );
DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1__9_), .Q(a_e_9_) );
DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_5__0_), .Q(b_e_0_) );
DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_5__1_), .Q(b_e_1_) );
DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_5__2_), .Q(b_e_2_) );
DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_5__3_), .Q(b_e_3_) );
DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_5__4_), .Q(b_e_4_) );
DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_5__5_), .Q(b_e_5_) );
DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_5__6_), .Q(b_e_6_) );
DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_5__7_), .Q(b_e_7_) );
DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_5__8_), .Q(b_e_8_) );
DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_5__9_), .Q(b_e_9_) );
DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_21__0_), .Q(z_e_0_) );
DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_21__1_), .Q(z_e_1_) );
DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21__2_), .Q(z_e_2_) );
DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_21__3_), .Q(z_e_3_) );
DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_21__4_), .Q(z_e_4_) );
DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_21__5_), .Q(z_e_5_) );
DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21__6_), .Q(z_e_6_) );
DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21__7_), .Q(z_e_7_) );
DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21__8_), .Q(z_e_8_) );
DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_21__9_), .Q(z_e_9_) );
DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3_), .Q(a_s) );
DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_7_), .Q(b_s) );
DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_23_), .Q(z_s) );
DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_11_), .Q(guard) );
DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_14_), .Q(round_bit) );
DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_19_), .Q(sticky) );
DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_12__0_), .Q(quotient_0_) );
DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_12__1_), .Q(quotient_1_) );
DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_12__2_), .Q(quotient_2_) );
DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__3_), .Q(quotient_3_) );
DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__4_), .Q(quotient_4_) );
DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__5_), .Q(quotient_5_) );
DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_12__6_), .Q(quotient_6_) );
DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__7_), .Q(quotient_7_) );
DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_12__8_), .Q(quotient_8_) );
DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__9_), .Q(quotient_9_) );
DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__10_), .Q(quotient_10_) );
DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12__11_), .Q(quotient_11_) );
DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__12_), .Q(quotient_12_) );
DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_12__13_), .Q(quotient_13_) );
DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__14_), .Q(quotient_14_) );
DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__15_), .Q(quotient_15_) );
DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__16_), .Q(quotient_16_) );
DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__17_), .Q(quotient_17_) );
DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__18_), .Q(quotient_18_) );
DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__19_), .Q(quotient_19_) );
DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__20_), .Q(quotient_20_) );
DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__21_), .Q(quotient_21_) );
DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__22_), .Q(quotient_22_) );
DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__23_), .Q(quotient_23_) );
DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12__24_), .Q(quotient_24_) );
DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12__25_), .Q(quotient_25_) );
DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_12__26_), .Q(quotient_26_) );
DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_10__0_), .Q(divisor_0_) );
DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_10__1_), .Q(divisor_1_) );
DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_10__2_), .Q(divisor_2_) );
DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__3_), .Q(divisor_3_) );
DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_10__4_), .Q(divisor_4_) );
DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__5_), .Q(divisor_5_) );
DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_10__6_), .Q(divisor_6_) );
DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__7_), .Q(divisor_7_) );
DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_10__8_), .Q(divisor_8_) );
DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__9_), .Q(divisor_9_) );
DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10__10_), .Q(divisor_10_) );
DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_10__11_), .Q(divisor_11_) );
DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_10__12_), .Q(divisor_12_) );
DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10__13_), .Q(divisor_13_) );
DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10__14_), .Q(divisor_14_) );
DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_10__15_), .Q(divisor_15_) );
DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_10__16_), .Q(divisor_16_) );
DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_10__17_), .Q(divisor_17_) );
DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__18_), .Q(divisor_18_) );
DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_10__19_), .Q(divisor_19_) );
DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__20_), .Q(divisor_20_) );
DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_10__21_), .Q(divisor_21_) );
DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_10__22_), .Q(divisor_22_) );
DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_10__23_), .Q(divisor_23_) );
DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__24_), .Q(divisor_24_) );
DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__25_), .Q(divisor_25_) );
DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__26_), .Q(divisor_26_) );
DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__27_), .Q(divisor_27_) );
DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_10__28_), .Q(divisor_28_) );
DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_10__29_), .Q(divisor_29_) );
DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_10__30_), .Q(divisor_30_) );
DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_10__31_), .Q(divisor_31_) );
DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__32_), .Q(divisor_32_) );
DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_10__33_), .Q(divisor_33_) );
DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_10__34_), .Q(divisor_34_) );
DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_10__35_), .Q(divisor_35_) );
DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_10__36_), .Q(divisor_36_) );
DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_10__37_), .Q(divisor_37_) );
DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__38_), .Q(divisor_38_) );
DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__39_), .Q(divisor_39_) );
DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_10__40_), .Q(divisor_40_) );
DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_10__41_), .Q(divisor_41_) );
DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_10__42_), .Q(divisor_42_) );
DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_10__43_), .Q(divisor_43_) );
DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_10__44_), .Q(divisor_44_) );
DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_10__45_), .Q(divisor_45_) );
DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_10__46_), .Q(divisor_46_) );
DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_10__47_), .Q(divisor_47_) );
DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_10__48_), .Q(divisor_48_) );
DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_10__49_), .Q(divisor_49_) );
DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_10__50_), .Q(divisor_50_) );
DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__0_), .Q(dividend_0_) );
DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__1_), .Q(dividend_1_) );
DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__2_), .Q(dividend_2_) );
DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__3_), .Q(dividend_3_) );
DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__4_), .Q(dividend_4_) );
DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__5_), .Q(dividend_5_) );
DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__6_), .Q(dividend_6_) );
DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__7_), .Q(dividend_7_) );
DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__8_), .Q(dividend_8_) );
DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__9_), .Q(dividend_9_) );
DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__10_), .Q(dividend_10_) );
DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__11_), .Q(dividend_11_) );
DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_9__12_), .Q(dividend_12_) );
DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_9__13_), .Q(dividend_13_) );
DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_9__14_), .Q(dividend_14_) );
DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__15_), .Q(dividend_15_) );
DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_9__16_), .Q(dividend_16_) );
DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__17_), .Q(dividend_17_) );
DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__18_), .Q(dividend_18_) );
DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__19_), .Q(dividend_19_) );
DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_9__20_), .Q(dividend_20_) );
DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__21_), .Q(dividend_21_) );
DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__22_), .Q(dividend_22_) );
DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__23_), .Q(dividend_23_) );
DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__24_), .Q(dividend_24_) );
DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__25_), .Q(dividend_25_) );
DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_9__26_), .Q(dividend_26_) );
DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_9__27_), .Q(dividend_27_) );
DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__28_), .Q(dividend_28_) );
DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__29_), .Q(dividend_29_) );
DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__30_), .Q(dividend_30_) );
DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_9__31_), .Q(dividend_31_) );
DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_9__32_), .Q(dividend_32_) );
DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__33_), .Q(dividend_33_) );
DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__34_), .Q(dividend_34_) );
DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__35_), .Q(dividend_35_) );
DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_9__36_), .Q(dividend_36_) );
DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__37_), .Q(dividend_37_) );
DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__38_), .Q(dividend_38_) );
DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_9__39_), .Q(dividend_39_) );
DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_9__40_), .Q(dividend_40_) );
DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_9__41_), .Q(dividend_41_) );
DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_9__42_), .Q(dividend_42_) );
DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_9__43_), .Q(dividend_43_) );
DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__44_), .Q(dividend_44_) );
DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__45_), .Q(dividend_45_) );
DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__46_), .Q(dividend_46_) );
DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_9__47_), .Q(dividend_47_) );
DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_9__48_), .Q(dividend_48_) );
DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_9__49_), .Q(dividend_49_) );
DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_9__50_), .Q(dividend_50_) );
DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__0_), .Q(remainder_0_) );
DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__1_), .Q(remainder_1_) );
DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__2_), .Q(remainder_2_) );
DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__3_), .Q(remainder_3_) );
DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__4_), .Q(remainder_4_) );
DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__5_), .Q(remainder_5_) );
DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__6_), .Q(remainder_6_) );
DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__7_), .Q(remainder_7_) );
DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__8_), .Q(remainder_8_) );
DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__9_), .Q(remainder_9_) );
DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13__10_), .Q(remainder_10_) );
DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13__11_), .Q(remainder_11_) );
DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_13__12_), .Q(remainder_12_) );
DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_13__13_), .Q(remainder_13_) );
DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_13__14_), .Q(remainder_14_) );
DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_13__15_), .Q(remainder_15_) );
DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13__16_), .Q(remainder_16_) );
DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13__17_), .Q(remainder_17_) );
DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13__18_), .Q(remainder_18_) );
DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_13__19_), .Q(remainder_19_) );
DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_13__20_), .Q(remainder_20_) );
DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_13__21_), .Q(remainder_21_) );
DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_13__22_), .Q(remainder_22_) );
DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_13__23_), .Q(remainder_23_) );
DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_13__24_), .Q(remainder_24_) );
DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_13__25_), .Q(remainder_25_) );
DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_13__26_), .Q(remainder_26_) );
DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_13__27_), .Q(remainder_27_) );
DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13__28_), .Q(remainder_28_) );
DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13__29_), .Q(remainder_29_) );
DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13__30_), .Q(remainder_30_) );
DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13__31_), .Q(remainder_31_) );
DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13__32_), .Q(remainder_32_) );
DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_13__33_), .Q(remainder_33_) );
DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_13__34_), .Q(remainder_34_) );
DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_13__35_), .Q(remainder_35_) );
DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_13__36_), .Q(remainder_36_) );
DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_13__37_), .Q(remainder_37_) );
DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_13__38_), .Q(remainder_38_) );
DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_13__39_), .Q(remainder_39_) );
DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_13__40_), .Q(remainder_40_) );
DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_13__41_), .Q(remainder_41_) );
DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_13__42_), .Q(remainder_42_) );
DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_13__43_), .Q(remainder_43_) );
DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13__44_), .Q(remainder_44_) );
DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_13__45_), .Q(remainder_45_) );
DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_13__46_), .Q(remainder_46_) );
DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_13__47_), .Q(remainder_47_) );
DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_13__48_), .Q(remainder_48_) );
DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_13__49_), .Q(remainder_49_) );
DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_13__50_), .Q(remainder_50_) );
DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8__0_), .Q(count_0_) );
DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8__1_), .Q(count_1_) );
DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8__2_), .Q(count_2_) );
DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8__3_), .Q(count_3_) );
DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8__4_), .Q(count_4_) );
DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_8__5_), .Q(count_5_) );
endmodule
