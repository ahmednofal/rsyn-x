module timer ( gnd, vdd, S_ADR_I, S_DAT_I, S_WE_I, S_STB_I, S_CYC_I, S_CTI_I, S_BTE_I, S_LOCK_I, S_SEL_I, CLK_I, RST_I, S_DAT_O, S_ACK_O, S_RTY_O, S_ERR_O, S_INT_O, RSTREQ_O, TOPULSE_O);

input gnd, vdd;
input S_WE_I;
input S_STB_I;
input S_CYC_I;
input S_LOCK_I;
input CLK_I;
input RST_I;
output S_ACK_O;
output S_RTY_O;
output S_ERR_O;
output S_INT_O;
output RSTREQ_O;
output TOPULSE_O;
input [31:0] S_ADR_I;
input [31:0] S_DAT_I;
input [2:0] S_CTI_I;
input [1:0] S_BTE_I;
input [3:0] S_SEL_I;
output [31:0] S_DAT_O;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_19__bF_buf4) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_19__bF_buf3) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_19__bF_buf2) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_19__bF_buf1) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_19__bF_buf0) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_86__bF_buf3) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_86__bF_buf2) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_86__bF_buf1) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_86__bF_buf0) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf7) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf6) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf5) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf4) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf3) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf2) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf1) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(RST_I), .Y(RST_I_bF_buf0) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf7) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf6) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf5) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf4) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf3) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf2) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf1) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(CLK_I), .Y(CLK_I_bF_buf0) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf5) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf4) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf3) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf2) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf1) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_58__bF_buf0) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(status_0_), .Y(status_0_bF_buf3) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(status_0_), .Y(status_0_bF_buf2) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(status_0_), .Y(status_0_bF_buf1) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(status_0_), .Y(status_0_bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_462__bF_buf4) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_462__bF_buf3) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_462__bF_buf2) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_462__bF_buf1) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_462__bF_buf0) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_469_), .Y(_510_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_15_), .B(_462__bF_buf1), .C(_510_), .Y(_511_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_511_), .Y(_528__15_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_58__bF_buf4), .C(_67_), .Y(_7__0_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_58__bF_buf4), .C(_99_), .Y(_7__1_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_58__bF_buf3), .C(_119_), .Y(_7__2_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_58__bF_buf0), .C(_140_), .Y(_7__3_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_58__bF_buf0), .C(_160_), .Y(_7__4_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_5_), .Y(_512_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_58__bF_buf5), .C(_178_), .Y(_7__5_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .Y(_513_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_58__bF_buf0), .C(_194_), .Y(_7__6_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_7_), .Y(_514_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_58__bF_buf3), .C(_214_), .Y(_7__7_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_58__bF_buf5), .C(_238_), .Y(_7__8_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_58__bF_buf5), .C(_276_), .Y(_7__9_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_58__bF_buf0), .C(_279_), .Y(_7__10_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_11_), .Y(_515_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_58__bF_buf0), .C(_304_), .Y(_7__11_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_58__bF_buf1), .C(_329_), .Y(_7__12_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_339_), .Y(_7__13_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_58__bF_buf2), .C(_373_), .Y(_7__14_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_58__bF_buf2), .C(_406_), .Y(_7__15_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(reg_wr), .B(dw04_cs), .Y(_516_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_2_), .B(_516_), .Y(_517_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(reg_stop), .C(latch_s_data_3_), .Y(_518_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_516_), .Y(_519_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_519_), .C(_518_), .Y(_10_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(status_2_), .Y(_520_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_18_), .C(reg_stop), .Y(_8_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(reg_ito), .Y(_521_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_0_), .B(_516_), .Y(_522_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_516_), .C(_522_), .Y(_6__0_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_1_), .B(_516_), .Y(_523_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_516_), .C(_523_), .Y(_6__1_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_521_), .Y(_524_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_0_), .B(_21_), .Y(_525_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(dw00_cs), .B(_525_), .C(_435_), .D(_524_), .Y(_11_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(s_ack_dly), .Y(_526_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(s_ack_2dly), .B(_526_), .Y(_527_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(reg_run), .B(_517_), .Y(_9_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_341_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_343_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_345_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_347_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_349_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_351_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_353_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_355_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_357_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_359_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_361_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_362_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_364_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_366_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_368_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_370_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_372_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_374_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_376_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_378_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_380_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_382_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_384_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_386_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_388_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_390_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_392_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_394_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_396_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_398_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_400_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_401_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_403_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_405_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_407_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_409_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_411_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_413_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_415_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_417_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_419_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_421_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_423_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_425_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_427_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_429_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_431_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_433_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_434_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_436_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_438_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_440_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_442_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_444_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf4), .Y(_446_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf0), .Y(_448_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_450_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf5), .Y(_452_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_454_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf1), .Y(_456_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf3), .Y(_458_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf7), .Y(_459_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_461_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf2), .Y(_463_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_465_) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(RSTREQ_O) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_527_), .Y(S_ACK_O) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_528__0_), .Y(S_DAT_O[0]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_528__1_), .Y(S_DAT_O[1]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_528__2_), .Y(S_DAT_O[2]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_528__3_), .Y(S_DAT_O[3]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_528__4_), .Y(S_DAT_O[4]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_528__5_), .Y(S_DAT_O[5]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_528__6_), .Y(S_DAT_O[6]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_528__7_), .Y(S_DAT_O[7]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_528__8_), .Y(S_DAT_O[8]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_528__9_), .Y(S_DAT_O[9]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_528__10_), .Y(S_DAT_O[10]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_528__11_), .Y(S_DAT_O[11]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_528__12_), .Y(S_DAT_O[12]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_528__13_), .Y(S_DAT_O[13]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_528__14_), .Y(S_DAT_O[14]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_528__15_), .Y(S_DAT_O[15]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[16]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[17]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[18]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[19]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[20]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[21]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[22]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[23]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[24]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[25]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[26]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[27]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[28]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[29]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[30]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_DAT_O[31]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_ERR_O) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_529_), .Y(S_INT_O) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(S_RTY_O) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_530_), .Y(TOPULSE_O) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(_16_), .Q(status_0_), .R(vdd), .S(_341_) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_15_), .Q(status_1_), .R(_343_), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_14_), .Q(status_2_), .R(_345_), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(_0_), .Q(_530_), .R(_347_), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(_7__0_), .Q(read_08_data_0_), .R(_349_), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_7__1_), .Q(read_08_data_1_), .R(_351_), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_7__2_), .Q(read_08_data_2_), .R(vdd), .S(_353_) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_7__3_), .Q(read_08_data_3_), .R(_355_), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_7__4_), .Q(read_08_data_4_), .R(vdd), .S(_357_) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_7__5_), .Q(read_08_data_5_), .R(_359_), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_7__6_), .Q(read_08_data_6_), .R(_361_), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_7__7_), .Q(read_08_data_7_), .R(_362_), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_7__8_), .Q(read_08_data_8_), .R(_364_), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_7__9_), .Q(read_08_data_9_), .R(_366_), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_7__10_), .Q(read_08_data_10_), .R(_368_), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_7__11_), .Q(read_08_data_11_), .R(_370_), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_7__12_), .Q(read_08_data_12_), .R(_372_), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_7__13_), .Q(read_08_data_13_), .R(_374_), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_7__14_), .Q(read_08_data_14_), .R(_376_), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_7__15_), .Q(read_08_data_15_), .R(_378_), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_10_), .Q(reg_stop), .R(_380_), .S(vdd) );
DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_8_), .Q(reg_run), .R(_382_), .S(vdd) );
DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_5__0_), .Q(internal_counter_0_), .R(_384_), .S(vdd) );
DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_5__1_), .Q(internal_counter_1_), .R(_386_), .S(vdd) );
DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_5__2_), .Q(internal_counter_2_), .R(_388_), .S(vdd) );
DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_5__3_), .Q(internal_counter_3_), .R(_390_), .S(vdd) );
DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_5__4_), .Q(internal_counter_4_), .R(_392_), .S(vdd) );
DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(_5__5_), .Q(internal_counter_5_), .R(_394_), .S(vdd) );
DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_5__6_), .Q(internal_counter_6_), .R(_396_), .S(vdd) );
DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_5__7_), .Q(internal_counter_7_), .R(_398_), .S(vdd) );
DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_5__8_), .Q(internal_counter_8_), .R(_400_), .S(vdd) );
DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_5__9_), .Q(internal_counter_9_), .R(_401_), .S(vdd) );
DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(_5__10_), .Q(internal_counter_10_), .R(_403_), .S(vdd) );
DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_5__11_), .Q(internal_counter_11_), .R(_405_), .S(vdd) );
DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_5__12_), .Q(internal_counter_12_), .R(_407_), .S(vdd) );
DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(_5__13_), .Q(internal_counter_13_), .R(_409_), .S(vdd) );
DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_5__14_), .Q(internal_counter_14_), .R(_411_), .S(vdd) );
DFFSR DFFSR_38 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_5__15_), .Q(internal_counter_15_), .R(_413_), .S(vdd) );
DFFSR DFFSR_39 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(s_ack_pre), .Q(s_ack_dly), .R(_415_), .S(vdd) );
DFFSR DFFSR_40 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(s_ack_dly), .Q(s_ack_2dly), .R(_417_), .S(vdd) );
DFFSR DFFSR_41 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(_13_), .Q(s_ack_pre), .R(_419_), .S(vdd) );
DFFSR DFFSR_42 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_6__0_), .Q(reg_ito), .R(_421_), .S(vdd) );
DFFSR DFFSR_43 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_6__1_), .Q(reg_cont), .R(_423_), .S(vdd) );
DFFSR DFFSR_44 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(_9_), .Q(reg_start), .R(_425_), .S(vdd) );
DFFSR DFFSR_45 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(_11_), .Q(_529_), .R(_427_), .S(vdd) );
DFFSR DFFSR_46 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_12_), .Q(reg_wr), .R(_429_), .S(vdd) );
DFFSR DFFSR_47 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(_1_), .Q(dw00_cs), .R(_431_), .S(vdd) );
DFFSR DFFSR_48 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_2_), .Q(dw04_cs), .R(_433_), .S(vdd) );
DFFSR DFFSR_49 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(_3_), .Q(dw08_cs), .R(_434_), .S(vdd) );
DFFSR DFFSR_50 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(_4_), .Q(dw0c_cs), .R(_436_), .S(vdd) );
DFFSR DFFSR_51 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf5), .D(S_DAT_I[0]), .Q(latch_s_data_0_), .R(_438_), .S(vdd) );
DFFSR DFFSR_52 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(S_DAT_I[1]), .Q(latch_s_data_1_), .R(_440_), .S(vdd) );
DFFSR DFFSR_53 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(S_DAT_I[2]), .Q(latch_s_data_2_), .R(_442_), .S(vdd) );
DFFSR DFFSR_54 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(S_DAT_I[3]), .Q(latch_s_data_3_), .R(_444_), .S(vdd) );
DFFSR DFFSR_55 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(S_DAT_I[4]), .Q(latch_s_data_4_), .R(_446_), .S(vdd) );
DFFSR DFFSR_56 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf6), .D(S_DAT_I[5]), .Q(latch_s_data_5_), .R(_448_), .S(vdd) );
DFFSR DFFSR_57 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(S_DAT_I[6]), .Q(latch_s_data_6_), .R(_450_), .S(vdd) );
DFFSR DFFSR_58 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf2), .D(S_DAT_I[7]), .Q(latch_s_data_7_), .R(_452_), .S(vdd) );
DFFSR DFFSR_59 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(S_DAT_I[8]), .Q(latch_s_data_8_), .R(_454_), .S(vdd) );
DFFSR DFFSR_60 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf3), .D(S_DAT_I[9]), .Q(latch_s_data_9_), .R(_456_), .S(vdd) );
DFFSR DFFSR_61 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf4), .D(S_DAT_I[10]), .Q(latch_s_data_10_), .R(_458_), .S(vdd) );
DFFSR DFFSR_62 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf7), .D(S_DAT_I[11]), .Q(latch_s_data_11_), .R(_459_), .S(vdd) );
DFFSR DFFSR_63 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(S_DAT_I[12]), .Q(latch_s_data_12_), .R(_461_), .S(vdd) );
DFFSR DFFSR_64 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(S_DAT_I[13]), .Q(latch_s_data_13_), .R(_463_), .S(vdd) );
DFFSR DFFSR_65 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf0), .D(S_DAT_I[14]), .Q(latch_s_data_14_), .R(_465_), .S(vdd) );
DFFSR DFFSR_66 ( .gnd(gnd), .vdd(vdd), .CLK(CLK_I_bF_buf1), .D(S_DAT_I[15]), .Q(latch_s_data_15_), .R(_17_), .S(vdd) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(RST_I_bF_buf6), .Y(_17_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(reg_start), .Y(_18_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(reg_stop), .B(_18_), .Y(_19_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(dw08_cs), .Y(_20_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(reg_wr), .Y(_21_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(status_0_bF_buf1), .Y(_22_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(_23_), .C(_19__bF_buf4), .Y(_24_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(reg_stop), .Y(_25_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_0_), .B(internal_counter_1_), .Y(_26_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_2_), .B(internal_counter_3_), .Y(_27_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .Y(_28_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_6_), .B(internal_counter_5_), .Y(_29_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_7_), .B(internal_counter_4_), .Y(_30_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .Y(_31_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_31_), .Y(_32_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_15_), .B(internal_counter_12_), .Y(_33_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_14_), .B(internal_counter_13_), .Y(_34_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .Y(_35_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_10_), .B(internal_counter_9_), .Y(_36_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_11_), .B(internal_counter_8_), .Y(_37_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .Y(_38_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_38_), .Y(_39_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_39_), .C(_25_), .Y(_40_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_39_), .Y(_41_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(reg_cont), .B(_41_), .C(status_2_), .Y(_42_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(_24_), .Y(_14_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(status_2_), .Y(_43_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .Y(_44_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .Y(_45_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .Y(_46_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .Y(_47_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .Y(_48_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_49_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49_), .C(reg_stop), .Y(_50_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .Y(_51_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_19__bF_buf2), .Y(_52_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_53_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_50_), .C(_53_), .Y(_15_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(reg_cont), .Y(_54_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49_), .Y(_55_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_55_), .Y(_56_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf4), .Y(_57_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_58_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_58__bF_buf3), .B(_57_), .C(status_0_bF_buf3), .Y(_59_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_56_), .C(_59_), .Y(_16_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[3]), .Y(_60_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[5]), .B(S_ADR_I[4]), .Y(_61_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .Y(_62_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[2]), .B(_62_), .Y(_1_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[2]), .Y(_63_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_62_), .Y(_2_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[3]), .B(_61_), .Y(_64_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(S_ADR_I[2]), .B(_64_), .Y(_3_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .Y(_4_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(S_STB_I), .B(S_CYC_I), .Y(_13_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(S_WE_I), .B(_13_), .Y(_65_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_12_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(reg_run), .B(_55_), .Y(_66_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_66_), .Y(_0_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_0_), .B(_58__bF_buf4), .Y(_67_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_0_), .Y(_69_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_10_), .B(read_08_data_11_), .Y(_70_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_8_), .B(read_08_data_9_), .Y(_71_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .Y(_72_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .B(read_08_data_1_), .Y(_73_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_2_), .B(read_08_data_3_), .Y(_74_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .Y(_75_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_4_), .B(read_08_data_5_), .Y(_76_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .B(read_08_data_7_), .Y(_77_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_78_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_75_), .C(_78_), .Y(_79_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_14_), .Y(_80_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_15_), .Y(_81_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .B(read_08_data_13_), .Y(_82_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_81_), .C(_82_), .Y(_83_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_79_), .C(_19__bF_buf3), .Y(_84_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .Y(_85_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_58__bF_buf3), .Y(_86_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_57_), .C(_86__bF_buf1), .Y(_87_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_69_), .C(_87_), .Y(_88_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_88_), .C(status_0_bF_buf3), .Y(_89_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(reg_stop), .B(_18_), .C(_58__bF_buf2), .Y(_90_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_91_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_91_), .Y(_92_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf1), .B(_67_), .Y(_93_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_92_), .C(status_1_), .Y(_94_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .B(_41_), .C(_69_), .Y(_95_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_58__bF_buf4), .B(_95_), .C(_67_), .Y(_96_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_69_), .C(_43_), .Y(_97_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_96_), .C(_97_), .Y(_98_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_89_), .C(_98_), .Y(_5__0_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_1_), .B(_58__bF_buf4), .Y(_99_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_1_), .Y(_101_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_1_), .Y(_102_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_102_), .Y(_103_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .B(read_08_data_1_), .C(_19__bF_buf1), .Y(_104_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_104_), .C(_86__bF_buf1), .Y(_105_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_101_), .C(_105_), .Y(_106_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_106_), .C(status_0_bF_buf3), .Y(_107_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(status_2_), .Y(_108_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_43_), .C(_108_), .Y(_109_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_1_), .B(_55_), .Y(_110_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_101_), .Y(_111_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_111_), .C(_41_), .Y(_112_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_112_), .C(_58__bF_buf3), .Y(_113_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_99_), .Y(_114_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_113_), .C(_109_), .Y(_115_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_91_), .Y(_116_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf1), .B(_99_), .Y(_117_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_116_), .C(status_1_), .Y(_118_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_107_), .C(_115_), .Y(_5__1_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_2_), .B(_58__bF_buf2), .Y(_119_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_2_), .Y(_121_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .B(read_08_data_1_), .C(read_08_data_2_), .Y(_122_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(_123_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_124_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_2_), .B(_124_), .C(_19__bF_buf1), .Y(_125_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_125_), .C(_86__bF_buf1), .Y(_126_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_121_), .C(_126_), .Y(_127_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_127_), .C(status_0_bF_buf3), .Y(_128_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_91_), .Y(_129_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf1), .B(_119_), .Y(_130_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_129_), .C(status_1_), .Y(_131_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_121_), .Y(_132_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49_), .C(_132_), .Y(_133_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_2_), .B(_32_), .C(_39_), .Y(_134_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_134_), .C(_58__bF_buf3), .Y(_135_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_2_), .Y(_136_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_86__bF_buf1), .C(_50_), .Y(_137_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_43_), .C(_108_), .Y(_138_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_137_), .C(_138_), .Y(_139_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_128_), .C(_139_), .Y(_5__2_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_3_), .B(_58__bF_buf4), .Y(_140_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_3_), .Y(_142_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_2_), .Y(_143_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_3_), .Y(_144_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_143_), .C(_144_), .Y(_145_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .Y(_146_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf2), .B(_146_), .Y(_147_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_147_), .C(_86__bF_buf2), .Y(_148_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_142_), .C(_148_), .Y(_149_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_149_), .C(status_0_bF_buf3), .Y(_150_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_121_), .C(_142_), .Y(_151_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_151_), .C(_86__bF_buf2), .Y(_152_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_144_), .C(_152_), .Y(_153_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_140_), .Y(_154_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_142_), .C(_43_), .Y(_155_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_153_), .C(_155_), .Y(_156_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_91_), .Y(_157_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf1), .B(_140_), .Y(_158_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_157_), .C(status_1_), .Y(_159_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_159_), .C(_150_), .Y(_5__3_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_4_), .B(_58__bF_buf4), .Y(_160_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_161_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_4_), .Y(_162_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_4_), .Y(_163_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_75_), .Y(_164_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_4_), .B(_146_), .C(_19__bF_buf2), .Y(_165_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_164_), .C(_86__bF_buf2), .Y(_166_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_162_), .C(_166_), .Y(_167_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_167_), .C(status_0_bF_buf0), .Y(_168_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_51_), .Y(_169_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_169_), .C(_52_), .D(_161_), .Y(_170_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_26_), .C(_27_), .Y(_171_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_4_), .B(_28_), .Y(_172_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_4_), .B(_41_), .C(_86__bF_buf2), .Y(_173_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_172_), .C(_173_), .Y(_174_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_160_), .Y(_175_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_43_), .C(_108_), .Y(_176_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_174_), .C(_176_), .Y(_177_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_168_), .C(_177_), .Y(_5__4_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_5_), .B(_58__bF_buf2), .Y(_178_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(_179_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_5_), .Y(_180_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_73_), .C(_74_), .Y(_181_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(read_08_data_5_), .Y(_182_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_5_), .B(_181_), .C(_19__bF_buf2), .Y(_183_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_86__bF_buf2), .Y(_184_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_180_), .C(_184_), .Y(_185_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_185_), .C(status_0_bF_buf0), .Y(_186_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_43_), .C(_108_), .Y(_187_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_180_), .Y(_188_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_5_), .B(_41_), .C(_86__bF_buf0), .Y(_189_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_189_), .C(_178_), .Y(_190_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_190_), .C(_187_), .Y(_191_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_51_), .Y(_192_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_192_), .C(_52_), .D(_179_), .Y(_193_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_186_), .C(_191_), .Y(_5__5_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_6_), .B(_58__bF_buf4), .Y(_194_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_195_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_6_), .Y(_196_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .C(_76_), .Y(_197_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(read_08_data_6_), .Y(_198_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .B(_197_), .C(_19__bF_buf2), .Y(_199_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_199_), .C(_86__bF_buf2), .Y(_200_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_196_), .C(_200_), .Y(_201_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_201_), .C(status_0_bF_buf0), .Y(_202_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_43_), .C(_108_), .Y(_203_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(_204_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_5_), .B(_171_), .C(internal_counter_6_), .Y(_205_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_204_), .C(_205_), .Y(_206_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .B(_41_), .C(_206_), .Y(_207_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_58__bF_buf0), .B(_207_), .C(_194_), .Y(_208_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_208_), .C(_203_), .Y(_209_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_91_), .Y(_210_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf2), .B(_194_), .Y(_211_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_210_), .C(status_1_), .Y(_212_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_202_), .C(_209_), .Y(_5__6_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf0), .Y(_213_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_7_), .B(_58__bF_buf3), .Y(_214_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_215_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_215_), .Y(_216_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .Y(_217_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_83_), .Y(_218_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_216_), .C(_57_), .Y(_219_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .B(_197_), .C(read_08_data_7_), .Y(_220_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_78_), .C(_57_), .Y(_221_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_220_), .C(_58__bF_buf5), .Y(_222_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_7_), .B(_219_), .C(_222_), .Y(_223_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_214_), .Y(_224_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_171_), .C(internal_counter_7_), .Y(_225_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_46_), .C(_225_), .Y(_226_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_226_), .Y(_227_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_7_), .B(_86__bF_buf0), .C(_55_), .Y(_228_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_229_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_40_), .Y(_230_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_230_), .Y(_231_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_7_), .Y(_232_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_232_), .C(_43_), .Y(_233_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_7_), .B(_86__bF_buf0), .C(_229_), .Y(_234_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_7_), .B(_19__bF_buf0), .Y(_235_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf0), .B(_234_), .C(_235_), .Y(_236_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(_236_), .C(_233_), .D(_231_), .Y(_237_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_224_), .C(_237_), .Y(_5__7_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_8_), .B(_58__bF_buf1), .Y(_238_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_8_), .B(_219_), .Y(_239_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_8_), .Y(_240_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_240_), .Y(_241_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_216_), .C(_19__bF_buf3), .Y(_242_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(_86__bF_buf3), .Y(_243_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_243_), .C(_238_), .Y(_244_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf2), .B(_244_), .Y(_245_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_8_), .Y(_246_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_91_), .Y(_247_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf4), .B(_238_), .Y(_248_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_247_), .C(status_1_), .Y(_249_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_31_), .C(_86__bF_buf0), .Y(_250_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_250_), .C(_246_), .Y(_251_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_58__bF_buf5), .Y(_252_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_32_), .C(_39_), .Y(_253_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_8_), .B(_28_), .C(_31_), .Y(_254_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .C(_58__bF_buf1), .Y(_255_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_8_), .B(_58__bF_buf1), .C(_254_), .D(_255_), .Y(_256_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_253_), .C(_40_), .Y(_257_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_257_), .C(status_2_), .Y(_258_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_258_), .C(_245_), .Y(_5__8_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_9_), .Y(_259_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_240_), .C(_259_), .Y(_260_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_75_), .C(_78_), .Y(_261_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf3), .B(_261_), .Y(_262_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_260_), .C(internal_counter_9_), .D(_219_), .Y(_263_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_263_), .Y(_264_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_9_), .Y(_265_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_58__bF_buf5), .Y(_266_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf1), .B(_266_), .C(_264_), .Y(_267_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_9_), .Y(_268_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_43_), .C(_108_), .Y(_269_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_268_), .C(_32_), .Y(_270_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_8_), .B(_46_), .C(internal_counter_9_), .Y(_271_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_9_), .B(_41_), .C(_86__bF_buf3), .Y(_272_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_271_), .C(_272_), .Y(_273_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_86__bF_buf3), .C(_50_), .Y(_274_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_273_), .C(_269_), .Y(_275_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_9_), .B(_58__bF_buf5), .Y(_276_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf3), .B(_276_), .C(_268_), .D(_91_), .Y(_277_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(_277_), .Y(_278_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_275_), .C(_267_), .Y(_5__9_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_10_), .B(_58__bF_buf0), .Y(_279_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_279_), .Y(_280_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_254_), .Y(_281_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49_), .C(_86__bF_buf1), .Y(_282_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_44_), .C(_45_), .Y(_283_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_9_), .B(_283_), .C(internal_counter_10_), .Y(_284_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(read_08_data_10_), .Y(_285_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_285_), .C(_281_), .D(_284_), .Y(_286_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_280_), .C(_286_), .Y(_287_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_10_), .B(_50_), .C(status_2_), .Y(_288_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_10_), .Y(_289_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_71_), .C(_216_), .Y(_290_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_10_), .B(_261_), .Y(_291_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf0), .B(_290_), .C(_291_), .Y(_292_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_10_), .Y(_293_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_293_), .C(_22_), .Y(_294_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf0), .B(_86__bF_buf0), .C(internal_counter_10_), .Y(_295_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf1), .B(_52_), .C(_280_), .Y(_296_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_295_), .C(_296_), .Y(_297_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_292_), .C(_297_), .Y(_298_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_287_), .C(_298_), .Y(_5__10_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_10_), .B(_270_), .C(internal_counter_11_), .Y(_299_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(_48_), .Y(_300_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_300_), .Y(_301_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_11_), .B(_35_), .C(_301_), .Y(_302_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_302_), .C(_58__bF_buf5), .Y(_303_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_11_), .B(_58__bF_buf3), .Y(_304_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_304_), .Y(_305_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_11_), .Y(_306_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_306_), .C(_43_), .Y(_307_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_303_), .C(_307_), .Y(_308_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(read_08_data_11_), .C(_57_), .Y(_309_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_11_), .B(_290_), .C(_309_), .Y(_310_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_306_), .C(_22_), .Y(_311_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf0), .B(_304_), .C(_306_), .D(_91_), .Y(_312_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(_312_), .Y(_313_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_304_), .C(_313_), .Y(_314_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_311_), .C(_314_), .Y(_315_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_308_), .Y(_5__11_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .B(_79_), .C(_19__bF_buf3), .Y(_316_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .Y(_317_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_72_), .C(_317_), .Y(_318_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_12_), .B(_219_), .C(_318_), .D(_316_), .Y(_319_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_86__bF_buf3), .B(_319_), .Y(_320_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_86__bF_buf3), .B(latch_s_data_12_), .Y(_321_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf2), .B(_321_), .C(_320_), .Y(_322_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_12_), .Y(_323_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_43_), .C(_108_), .Y(_324_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_323_), .Y(_325_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .B(_41_), .C(_86__bF_buf3), .Y(_326_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_12_), .B(_58__bF_buf1), .C(_40_), .Y(_327_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_325_), .C(_327_), .Y(_328_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_12_), .B(_58__bF_buf1), .Y(_329_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf4), .B(_329_), .C(_323_), .D(_91_), .Y(_330_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(status_1_), .B(_330_), .C(_324_), .D(_328_), .Y(_331_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_322_), .Y(_5__12_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_13_), .Y(_332_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_43_), .C(_108_), .Y(_333_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_12_), .B(_300_), .Y(_334_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_334_), .Y(_335_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_12_), .B(_300_), .C(internal_counter_13_), .Y(_336_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(read_08_data_13_), .Y(_337_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_337_), .C(_336_), .D(_335_), .Y(_338_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_13_), .B(_58__bF_buf2), .Y(_339_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_339_), .Y(_340_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_338_), .C(_333_), .Y(_342_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_82_), .C(_216_), .Y(_344_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .B(_79_), .C(read_08_data_13_), .Y(_346_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf3), .B(_344_), .C(_346_), .Y(_348_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_332_), .C(_22_), .Y(_350_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_13_), .B(status_1_), .Y(_352_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_339_), .Y(_354_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf1), .B(_52_), .C(_354_), .Y(_356_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_352_), .C(_356_), .Y(_358_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_348_), .C(_358_), .Y(_360_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_342_), .Y(_5__13_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_48_), .C(_32_), .Y(_363_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_13_), .B(_363_), .C(internal_counter_14_), .Y(_365_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_334_), .Y(_367_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(read_08_data_14_), .Y(_369_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_369_), .C(_365_), .D(_367_), .Y(_371_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_14_), .B(_58__bF_buf2), .Y(_373_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_55_), .C(_373_), .Y(_375_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_14_), .Y(_377_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_377_), .C(_43_), .Y(_379_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_371_), .C(_379_), .Y(_381_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_80_), .Y(_383_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_344_), .Y(_385_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_383_), .C(_19__bF_buf4), .Y(_387_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_377_), .C(_22_), .Y(_389_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_14_), .B(status_1_), .Y(_391_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_373_), .Y(_393_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf2), .B(_52_), .C(_393_), .Y(_395_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_391_), .C(_395_), .Y(_397_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .C(_397_), .Y(_399_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_399_), .Y(_5__14_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(internal_counter_15_), .Y(_402_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_34_), .C(_402_), .Y(_404_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(latch_s_data_15_), .B(_58__bF_buf2), .Y(_406_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_58__bF_buf1), .Y(_408_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_32_), .C(_39_), .Y(_410_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_410_), .C(_50_), .Y(_412_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_15_), .Y(_414_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_414_), .C(_43_), .Y(_416_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_404_), .C(_416_), .Y(_418_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_15_), .B(_84_), .Y(_420_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_14_), .B(_344_), .C(read_08_data_15_), .Y(_422_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_422_), .C(_420_), .Y(_424_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_424_), .Y(_426_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_406_), .Y(_428_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_19__bF_buf4), .B(_406_), .C(_414_), .D(_91_), .Y(_430_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(status_0_bF_buf2), .B(_428_), .C(status_1_), .D(_430_), .Y(_432_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_432_), .C(_426_), .Y(_5__15_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_529_), .Y(_435_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(S_STB_I), .Y(_437_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(S_WE_I), .B(_437_), .Y(_439_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(dw00_cs), .B(_439_), .Y(_441_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_439_), .Y(_443_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_443_), .Y(_445_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(dw04_cs), .B(_439_), .Y(_447_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(dw0c_cs), .B(_439_), .Y(_449_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(internal_counter_0_), .B(_20_), .Y(_451_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_449_), .C(_447_), .Y(_453_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_0_), .B(_445_), .C(_453_), .Y(_455_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(reg_ito), .B(_447_), .C(_441_), .Y(_457_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_441_), .C(_457_), .D(_455_), .Y(_528__0_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(reg_run), .Y(_460_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(_445_), .Y(_462_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_449_), .Y(_464_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_462__bF_buf3), .C(_447_), .Y(_466_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_462__bF_buf3), .C(_466_), .Y(_467_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(reg_cont), .B(_447_), .C(_441_), .Y(_468_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_441_), .C(_468_), .D(_467_), .Y(_528__1_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(dw04_cs), .B(dw00_cs), .C(_439_), .Y(_469_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_449_), .C(_462__bF_buf3), .Y(_470_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_469_), .Y(_471_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_2_), .B(_462__bF_buf4), .C(_471_), .Y(_472_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_472_), .Y(_528__2_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_449_), .C(_462__bF_buf2), .Y(_473_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_469_), .Y(_474_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_3_), .B(_462__bF_buf2), .C(_474_), .Y(_475_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_475_), .Y(_528__3_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_449_), .C(_462__bF_buf2), .Y(_476_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_469_), .Y(_477_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_4_), .B(_462__bF_buf2), .C(_477_), .Y(_478_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_478_), .Y(_528__4_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_449_), .C(_462__bF_buf4), .Y(_479_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_469_), .Y(_480_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_5_), .B(_462__bF_buf4), .C(_480_), .Y(_481_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_481_), .Y(_528__5_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_449_), .C(_462__bF_buf4), .Y(_482_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_469_), .Y(_483_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_6_), .B(_462__bF_buf2), .C(_483_), .Y(_484_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_484_), .Y(_528__6_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_449_), .C(_462__bF_buf4), .Y(_485_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_469_), .Y(_486_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_7_), .B(_462__bF_buf2), .C(_486_), .Y(_487_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_487_), .Y(_528__7_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_449_), .C(_462__bF_buf1), .Y(_488_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_469_), .Y(_489_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_8_), .B(_462__bF_buf1), .C(_489_), .Y(_490_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_528__8_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_449_), .C(_462__bF_buf1), .Y(_491_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_469_), .Y(_492_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_9_), .B(_462__bF_buf0), .C(_492_), .Y(_493_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_493_), .Y(_528__9_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_449_), .C(_462__bF_buf0), .Y(_494_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_469_), .Y(_495_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_10_), .B(_462__bF_buf4), .C(_495_), .Y(_496_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_496_), .Y(_528__10_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_449_), .C(_462__bF_buf0), .Y(_497_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_469_), .Y(_498_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_11_), .B(_462__bF_buf0), .C(_498_), .Y(_499_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_499_), .Y(_528__11_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_449_), .C(_462__bF_buf1), .Y(_500_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_469_), .Y(_501_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_12_), .B(_462__bF_buf1), .C(_501_), .Y(_502_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_502_), .Y(_528__12_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_449_), .C(_462__bF_buf0), .Y(_503_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_469_), .Y(_504_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_13_), .B(_462__bF_buf0), .C(_504_), .Y(_505_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_505_), .Y(_528__13_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_449_), .C(_462__bF_buf3), .Y(_506_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_469_), .Y(_507_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(read_08_data_14_), .B(_462__bF_buf3), .C(_507_), .Y(_508_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_508_), .Y(_528__14_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_449_), .C(_462__bF_buf3), .Y(_509_) );
endmodule
