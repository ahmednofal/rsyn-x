magic
tech scmos
magscale 1 2
timestamp 1522732896
<< metal1 >>
rect 3112 4606 3113 4614
rect 3121 4606 3123 4614
rect 3131 4606 3133 4614
rect 3141 4606 3143 4614
rect 3151 4606 3160 4614
rect 4653 4557 4700 4563
rect 5796 4556 5804 4564
rect 6068 4557 6083 4563
rect 332 4537 371 4543
rect 1357 4537 1372 4543
rect 1588 4537 1612 4543
rect 1620 4537 1635 4543
rect 1812 4537 1827 4543
rect 3405 4537 3420 4543
rect 3868 4537 3892 4543
rect 4093 4543 4099 4556
rect 4093 4537 4115 4543
rect 4148 4537 4163 4543
rect 4765 4537 4780 4543
rect 5485 4537 5523 4543
rect 5821 4537 5859 4543
rect 6100 4537 6131 4543
rect 93 4517 131 4523
rect 260 4517 275 4523
rect 676 4517 707 4523
rect 1268 4517 1283 4523
rect 1636 4517 1651 4523
rect 1748 4517 1763 4523
rect 1773 4517 1788 4523
rect 1853 4517 1875 4523
rect 2173 4517 2204 4523
rect 2308 4517 2323 4523
rect 2349 4517 2387 4523
rect 29 4497 67 4503
rect 84 4496 92 4504
rect 653 4497 691 4503
rect 1005 4497 1020 4503
rect 1652 4496 1660 4504
rect 2324 4496 2332 4504
rect 2349 4497 2355 4517
rect 2701 4517 2739 4523
rect 2733 4497 2739 4517
rect 3268 4517 3283 4523
rect 3405 4517 3443 4523
rect 3405 4497 3411 4517
rect 3949 4517 3964 4523
rect 4125 4517 4163 4523
rect 4189 4517 4204 4523
rect 4157 4497 4163 4517
rect 4548 4517 4563 4523
rect 4765 4517 4803 4523
rect 4765 4497 4771 4517
rect 5332 4517 5347 4523
rect 5565 4517 5580 4523
rect 5940 4517 5971 4523
rect 5412 4496 5420 4504
rect 5716 4497 5731 4503
rect 3661 4477 3676 4483
rect 4868 4476 4874 4484
rect 6020 4476 6022 4484
rect 6269 4477 6300 4483
rect 1576 4406 1577 4414
rect 1585 4406 1587 4414
rect 1595 4406 1597 4414
rect 1605 4406 1607 4414
rect 1615 4406 1624 4414
rect 4664 4406 4665 4414
rect 4673 4406 4675 4414
rect 4683 4406 4685 4414
rect 4693 4406 4695 4414
rect 4703 4406 4712 4414
rect 970 4376 972 4384
rect 2282 4376 2284 4384
rect 2810 4376 2812 4384
rect 2954 4376 2956 4384
rect 3530 4376 3532 4384
rect 5786 4376 5788 4384
rect 6154 4376 6156 4384
rect 5914 4356 5916 4364
rect 1034 4336 1036 4344
rect 2189 4337 2204 4343
rect 2621 4337 2636 4343
rect 3341 4337 3356 4343
rect 5636 4336 5638 4344
rect 269 4297 300 4303
rect 461 4297 476 4303
rect 740 4297 755 4303
rect 973 4297 1004 4303
rect 1117 4297 1139 4303
rect 1245 4297 1260 4303
rect 1780 4297 1811 4303
rect 1901 4297 1916 4303
rect 2077 4297 2092 4303
rect 2253 4303 2259 4323
rect 2221 4297 2259 4303
rect 2509 4297 2540 4303
rect 3453 4297 3500 4303
rect 3629 4303 3635 4323
rect 3629 4297 3667 4303
rect 4525 4303 4531 4323
rect 4637 4317 4652 4323
rect 4493 4297 4531 4303
rect 5181 4303 5187 4323
rect 5149 4297 5187 4303
rect 5213 4297 5228 4303
rect 5588 4297 5603 4303
rect 5668 4297 5715 4303
rect 5725 4297 5756 4303
rect 6109 4297 6147 4303
rect 6157 4297 6172 4303
rect 188 4277 212 4283
rect 1053 4277 1068 4283
rect 1469 4277 1484 4283
rect 1469 4257 1475 4277
rect 1924 4277 1939 4283
rect 2333 4277 2355 4283
rect 2436 4277 2452 4283
rect 3069 4277 3091 4283
rect 3677 4277 3692 4283
rect 3709 4277 3731 4283
rect 4212 4277 4227 4283
rect 4237 4277 4252 4283
rect 4468 4277 4483 4283
rect 4573 4277 4588 4283
rect 4660 4277 4723 4283
rect 5965 4277 5980 4283
rect 6068 4277 6083 4283
rect 6228 4277 6243 4283
rect 3101 4257 3116 4263
rect 3428 4256 3430 4264
rect 3693 4257 3699 4276
rect 4637 4257 4652 4263
rect 5988 4257 6003 4263
rect 6052 4257 6067 4263
rect 6253 4257 6268 4263
rect 2420 4236 2422 4244
rect 3050 4236 3052 4244
rect 3748 4236 3750 4244
rect 3978 4236 3980 4244
rect 5284 4236 5288 4244
rect 3112 4206 3113 4214
rect 3121 4206 3123 4214
rect 3131 4206 3133 4214
rect 3141 4206 3143 4214
rect 3151 4206 3160 4214
rect 1370 4176 1372 4184
rect 2936 4176 2940 4184
rect 3636 4176 3638 4184
rect 3992 4176 3996 4184
rect 6084 4176 6086 4184
rect 1604 4157 1651 4163
rect 3156 4157 3203 4163
rect 253 4137 275 4143
rect 1149 4137 1171 4143
rect 1309 4137 1324 4143
rect 1917 4137 1932 4143
rect 1997 4137 2019 4143
rect 2220 4137 2259 4143
rect 2509 4137 2531 4143
rect 2541 4137 2556 4143
rect 292 4117 307 4123
rect 916 4117 931 4123
rect 980 4117 995 4123
rect 1069 4117 1107 4123
rect 1133 4117 1148 4123
rect 996 4096 1004 4104
rect 1101 4097 1107 4117
rect 1293 4117 1308 4123
rect 1604 4117 1644 4123
rect 1284 4096 1292 4104
rect 1972 4096 1980 4104
rect 2493 4084 2499 4136
rect 3572 4117 3587 4123
rect 3773 4117 3779 4176
rect 4637 4157 4684 4163
rect 5444 4157 5459 4163
rect 4444 4144 4452 4148
rect 5933 4144 5939 4163
rect 4788 4137 4803 4143
rect 5069 4137 5084 4143
rect 5133 4137 5171 4143
rect 5524 4137 5539 4143
rect 5549 4124 5555 4143
rect 5796 4137 5811 4143
rect 5965 4137 6003 4143
rect 6068 4137 6083 4143
rect 6109 4137 6124 4143
rect 4100 4117 4115 4123
rect 4532 4117 4547 4123
rect 5028 4117 5043 4123
rect 5277 4117 5315 4123
rect 4141 4097 4156 4103
rect 5277 4097 5283 4117
rect 5508 4117 5523 4123
rect 5316 4096 5324 4104
rect 5517 4097 5523 4117
rect 5556 4117 5619 4123
rect 5684 4117 5699 4123
rect 5725 4117 5763 4123
rect 5725 4097 5731 4117
rect 5780 4117 5827 4123
rect 5837 4117 5875 4123
rect 5901 4117 5916 4123
rect 5869 4097 5875 4117
rect 6132 4117 6140 4123
rect 6173 4117 6188 4123
rect 6164 4096 6172 4104
rect 6205 4097 6220 4103
rect 314 4076 316 4084
rect 2628 4077 2643 4083
rect 2676 4077 2723 4083
rect 372 4056 374 4064
rect 2717 4057 2723 4077
rect 2964 4077 2995 4083
rect 1796 4036 1798 4044
rect 3156 4037 3180 4043
rect 5188 4036 5190 4044
rect 5898 4036 5900 4044
rect 1576 4006 1577 4014
rect 1585 4006 1587 4014
rect 1595 4006 1597 4014
rect 1605 4006 1607 4014
rect 1615 4006 1624 4014
rect 4664 4006 4665 4014
rect 4673 4006 4675 4014
rect 4683 4006 4685 4014
rect 4693 4006 4695 4014
rect 4703 4006 4712 4014
rect 180 3976 182 3984
rect 490 3976 492 3984
rect 1364 3976 1366 3984
rect 1802 3976 1804 3984
rect 5956 3976 5958 3984
rect 797 3937 812 3943
rect 4045 3937 4076 3943
rect 420 3916 428 3924
rect 868 3916 876 3924
rect 205 3897 259 3903
rect 893 3903 899 3923
rect 1108 3916 1116 3924
rect 2701 3917 2716 3923
rect 3117 3917 3164 3923
rect 893 3897 931 3903
rect 1005 3897 1020 3903
rect 1140 3897 1148 3903
rect 1828 3897 1843 3903
rect 557 3877 572 3883
rect 829 3877 844 3883
rect 989 3877 1036 3883
rect 1156 3877 1171 3883
rect 1501 3877 1516 3883
rect 1837 3877 1843 3897
rect 2573 3897 2596 3903
rect 2588 3892 2596 3897
rect 2868 3897 2883 3903
rect 3117 3903 3123 3917
rect 3101 3897 3123 3903
rect 2013 3877 2035 3883
rect 2077 3877 2092 3883
rect 2996 3877 3011 3883
rect 3085 3877 3148 3883
rect 3853 3877 3875 3883
rect 4045 3877 4051 3937
rect 5028 3937 5043 3943
rect 5770 3936 5772 3944
rect 4077 3897 4083 3916
rect 4132 3897 4147 3903
rect 4333 3903 4339 3923
rect 5412 3916 5420 3924
rect 6237 3917 6252 3923
rect 4292 3897 4307 3903
rect 4333 3897 4371 3903
rect 5101 3897 5155 3903
rect 5261 3897 5283 3903
rect 5661 3903 5667 3916
rect 5549 3897 5571 3903
rect 5661 3897 5699 3903
rect 5796 3897 5811 3903
rect 5924 3897 5955 3903
rect 6221 3897 6236 3903
rect 4333 3877 4348 3883
rect 4381 3877 4404 3883
rect 4396 3872 4404 3877
rect 5060 3877 5075 3883
rect 5204 3877 5219 3883
rect 5229 3877 5267 3883
rect 29 3857 44 3863
rect 1261 3857 1283 3863
rect 1453 3857 1475 3863
rect 1693 3857 1715 3863
rect 1885 3857 1907 3863
rect 4020 3856 4028 3864
rect 4668 3863 4676 3872
rect 4668 3857 4700 3863
rect 5229 3857 5235 3877
rect 5380 3877 5395 3883
rect 5844 3877 5859 3883
rect 6109 3877 6140 3883
rect 5636 3856 5644 3864
rect 2740 3836 2742 3844
rect 3576 3836 3580 3844
rect 3780 3837 3795 3843
rect 3834 3836 3836 3844
rect 3112 3806 3113 3814
rect 3121 3806 3123 3814
rect 3131 3806 3133 3814
rect 3141 3806 3143 3814
rect 3151 3806 3160 3814
rect 164 3776 166 3784
rect 468 3776 470 3784
rect 1492 3776 1494 3784
rect 1572 3776 1574 3784
rect 1908 3776 1910 3784
rect 2794 3776 2796 3784
rect 3796 3776 3798 3784
rect 4701 3777 4723 3783
rect 221 3737 259 3743
rect 392 3737 412 3743
rect 452 3737 460 3743
rect 556 3743 564 3744
rect 548 3737 564 3743
rect 884 3737 899 3743
rect 1124 3737 1139 3743
rect 1453 3743 1459 3763
rect 1725 3757 1747 3763
rect 4701 3763 4707 3777
rect 4996 3776 4998 3784
rect 4653 3757 4707 3763
rect 1453 3737 1468 3743
rect 1773 3737 1804 3743
rect 1892 3737 1907 3743
rect 2093 3737 2115 3743
rect 109 3717 140 3723
rect 180 3717 195 3723
rect 596 3717 611 3723
rect 973 3717 988 3723
rect 1197 3717 1212 3723
rect 1332 3717 1347 3723
rect 1613 3717 1660 3723
rect 1732 3717 1747 3723
rect 2036 3717 2051 3723
rect 2109 3723 2115 3737
rect 2132 3737 2147 3743
rect 3757 3737 3779 3743
rect 3876 3737 3891 3743
rect 4308 3737 4323 3743
rect 5108 3737 5123 3743
rect 5309 3737 5331 3743
rect 5540 3737 5560 3743
rect 5709 3737 5724 3743
rect 5764 3737 5772 3743
rect 5805 3737 5820 3743
rect 6196 3737 6211 3743
rect 6221 3737 6252 3743
rect 2109 3717 2131 3723
rect 2237 3717 2252 3723
rect 125 3697 140 3703
rect 420 3697 435 3703
rect 2125 3697 2131 3717
rect 2749 3717 2764 3723
rect 2781 3697 2787 3736
rect 3117 3717 3196 3723
rect 3348 3717 3356 3723
rect 3501 3717 3516 3723
rect 3645 3717 3683 3723
rect 2820 3697 2835 3703
rect 3172 3697 3203 3703
rect 3220 3696 3228 3704
rect 3677 3697 3683 3717
rect 4285 3717 4300 3723
rect 5396 3717 5411 3723
rect 5588 3717 5603 3723
rect 5613 3717 5651 3723
rect 3988 3677 4003 3683
rect 298 3656 300 3664
rect 3997 3657 4003 3677
rect 5693 3677 5724 3683
rect 970 3636 972 3644
rect 4676 3637 4700 3643
rect 1576 3606 1577 3614
rect 1585 3606 1587 3614
rect 1595 3606 1597 3614
rect 1605 3606 1607 3614
rect 1615 3606 1624 3614
rect 4664 3606 4665 3614
rect 4673 3606 4675 3614
rect 4683 3606 4685 3614
rect 4693 3606 4695 3614
rect 4703 3606 4712 3614
rect 500 3576 502 3584
rect 2154 3576 2156 3584
rect 3002 3576 3004 3584
rect 3082 3576 3084 3584
rect 3322 3576 3324 3584
rect 5226 3576 5228 3584
rect 5588 3576 5590 3584
rect 5764 3576 5766 3584
rect 5988 3576 5990 3584
rect 2436 3556 2438 3564
rect 893 3537 908 3543
rect 1476 3537 1507 3543
rect 2842 3536 2844 3544
rect 3748 3537 3779 3543
rect 4340 3537 4355 3543
rect 4740 3537 4755 3543
rect 580 3517 595 3523
rect 1252 3516 1260 3524
rect 1604 3517 1635 3523
rect 1757 3517 1779 3523
rect 84 3497 99 3503
rect 109 3497 124 3503
rect 1044 3497 1059 3503
rect 1236 3497 1251 3503
rect 1389 3497 1420 3503
rect 1629 3503 1635 3517
rect 1924 3516 1932 3524
rect 3732 3517 3747 3523
rect 3949 3517 3964 3523
rect 4541 3517 4556 3523
rect 1629 3497 1651 3503
rect 3325 3497 3340 3503
rect 3860 3497 3875 3503
rect 4285 3497 4300 3503
rect 4564 3497 4579 3503
rect 4829 3503 4835 3523
rect 4829 3497 4867 3503
rect 4980 3497 5011 3503
rect 5124 3497 5155 3503
rect 5357 3497 5379 3503
rect 5613 3503 5619 3523
rect 5572 3497 5587 3503
rect 5613 3497 5651 3503
rect 5789 3503 5795 3523
rect 6013 3517 6035 3523
rect 5709 3497 5763 3503
rect 5789 3497 5827 3503
rect 5949 3497 5987 3503
rect 6084 3497 6099 3503
rect 6196 3497 6227 3503
rect 28 3477 44 3483
rect 28 3476 36 3477
rect 125 3477 140 3483
rect 957 3477 972 3483
rect 1085 3477 1123 3483
rect 1117 3464 1123 3477
rect 1325 3477 1363 3483
rect 1604 3477 1644 3483
rect 1821 3477 1836 3483
rect 1997 3477 2028 3483
rect 2180 3477 2195 3483
rect 2621 3477 2627 3496
rect 3100 3492 3108 3496
rect 3108 3477 3164 3483
rect 3405 3477 3420 3483
rect 4829 3477 4844 3483
rect 4877 3477 4900 3483
rect 1757 3457 1763 3476
rect 2236 3472 2244 3476
rect 4892 3472 4900 3477
rect 5309 3477 5324 3483
rect 5428 3477 5443 3483
rect 6084 3477 6115 3483
rect 3156 3457 3171 3463
rect 237 3437 268 3443
rect 3693 3437 3708 3443
rect 4052 3436 4056 3444
rect 3112 3406 3113 3414
rect 3121 3406 3123 3414
rect 3131 3406 3133 3414
rect 3141 3406 3143 3414
rect 3151 3406 3160 3414
rect 1492 3376 1494 3384
rect 3140 3377 3164 3383
rect 3594 3376 3596 3384
rect 660 3356 668 3364
rect 1428 3356 1436 3364
rect 845 3337 883 3343
rect 973 3337 1011 3343
rect 973 3324 979 3337
rect 1284 3337 1315 3343
rect 1565 3337 1612 3343
rect 1668 3337 1683 3343
rect 620 3317 636 3323
rect 620 3312 628 3317
rect 701 3317 716 3323
rect 1549 3317 1651 3323
rect 1677 3317 1683 3337
rect 1869 3337 1884 3343
rect 2141 3337 2156 3343
rect 2356 3337 2364 3343
rect 2461 3343 2467 3363
rect 3757 3357 3772 3363
rect 2461 3337 2476 3343
rect 2205 3317 2211 3336
rect 2509 3324 2515 3343
rect 2253 3317 2300 3323
rect 2685 3323 2691 3343
rect 2861 3337 2876 3343
rect 3085 3337 3100 3343
rect 3540 3337 3548 3343
rect 2685 3317 2700 3323
rect 3309 3317 3356 3323
rect 3396 3317 3427 3323
rect 3437 3317 3475 3323
rect 3517 3317 3532 3323
rect 852 3297 867 3303
rect 1396 3297 1411 3303
rect 2052 3296 2060 3304
rect 2244 3296 2252 3304
rect 2836 3296 2844 3304
rect 3693 3284 3699 3343
rect 3780 3337 3795 3343
rect 3709 3317 3740 3323
rect 3789 3317 3795 3337
rect 4068 3337 4083 3343
rect 4221 3343 4227 3363
rect 4756 3357 4771 3363
rect 4221 3337 4236 3343
rect 4765 3343 4771 3357
rect 4765 3337 4787 3343
rect 4829 3337 4844 3343
rect 4892 3343 4900 3348
rect 4877 3337 4900 3343
rect 5124 3337 5139 3343
rect 5341 3337 5363 3343
rect 5677 3337 5699 3343
rect 5764 3337 5779 3343
rect 5789 3337 5827 3343
rect 5853 3343 5859 3363
rect 5844 3337 5859 3343
rect 6148 3337 6163 3343
rect 6189 3337 6243 3343
rect 3933 3317 3964 3323
rect 4253 3317 4291 3323
rect 4285 3297 4291 3317
rect 4436 3317 4467 3323
rect 4628 3317 4659 3323
rect 4829 3317 4867 3323
rect 4308 3296 4316 3304
rect 4829 3297 4835 3317
rect 5101 3317 5139 3323
rect 5133 3297 5139 3317
rect 5277 3317 5308 3323
rect 5277 3297 5283 3317
rect 5444 3317 5459 3323
rect 5492 3317 5523 3323
rect 5604 3317 5651 3323
rect 5725 3317 5763 3323
rect 5485 3297 5500 3303
rect 5757 3297 5763 3317
rect 5860 3317 5875 3323
rect 2572 3277 2595 3283
rect 2909 3277 2932 3283
rect 2730 3236 2732 3244
rect 2788 3236 2790 3244
rect 3044 3236 3046 3244
rect 5908 3236 5910 3244
rect 1576 3206 1577 3214
rect 1585 3206 1587 3214
rect 1595 3206 1597 3214
rect 1605 3206 1607 3214
rect 1615 3206 1624 3214
rect 4664 3206 4665 3214
rect 4673 3206 4675 3214
rect 4683 3206 4685 3214
rect 4693 3206 4695 3214
rect 4703 3206 4712 3214
rect 1834 3176 1836 3184
rect 1930 3176 1932 3184
rect 2330 3176 2332 3184
rect 3348 3176 3350 3184
rect 5844 3176 5846 3184
rect 1588 3157 1612 3163
rect 1469 3137 1484 3143
rect 2858 3136 2860 3144
rect 3796 3136 3798 3144
rect 3988 3136 3992 3144
rect 4532 3137 4547 3143
rect 4804 3136 4806 3144
rect 5581 3137 5596 3143
rect 5914 3136 5916 3144
rect 228 3116 236 3124
rect 397 3117 412 3123
rect 1652 3116 1660 3124
rect 77 3097 92 3103
rect 292 3097 307 3103
rect 1517 3097 1532 3103
rect 1517 3084 1523 3097
rect 1572 3097 1644 3103
rect 1677 3103 1683 3123
rect 2436 3116 2444 3124
rect 3140 3117 3155 3123
rect 1677 3097 1715 3103
rect 2397 3097 2412 3103
rect 1028 3077 1043 3083
rect 1092 3077 1107 3083
rect 1208 3076 1212 3084
rect 1572 3077 1628 3083
rect 2013 3077 2028 3083
rect 477 3057 508 3063
rect 868 3056 876 3064
rect 1000 3057 1027 3063
rect 2013 3057 2019 3077
rect 2173 3077 2188 3083
rect 2221 3077 2259 3083
rect 2397 3077 2403 3097
rect 2708 3097 2723 3103
rect 3149 3103 3155 3117
rect 3149 3097 3203 3103
rect 3332 3097 3347 3103
rect 3540 3097 3571 3103
rect 3652 3097 3667 3103
rect 3757 3097 3795 3103
rect 4045 3097 4076 3103
rect 2749 3077 2764 3083
rect 3421 3077 3436 3083
rect 3693 3077 3708 3083
rect 2372 3056 2380 3064
rect 3156 3057 3203 3063
rect 3693 3057 3699 3077
rect 4045 3077 4051 3097
rect 4157 3097 4195 3103
rect 4829 3103 4835 3123
rect 5444 3116 5452 3124
rect 4788 3097 4803 3103
rect 4829 3097 4867 3103
rect 5284 3097 5299 3103
rect 5309 3097 5324 3103
rect 5357 3097 5379 3103
rect 5389 3097 5420 3103
rect 5476 3097 5491 3103
rect 5773 3097 5788 3103
rect 5869 3103 5875 3123
rect 5988 3117 6003 3123
rect 6013 3117 6051 3123
rect 6244 3116 6252 3124
rect 6269 3117 6284 3123
rect 5869 3097 5907 3103
rect 6141 3097 6156 3103
rect 6196 3097 6243 3103
rect 4772 3077 4787 3083
rect 5492 3077 5507 3083
rect 5613 3077 5651 3083
rect 5805 3077 5827 3083
rect 3812 3057 3836 3063
rect 5380 3057 5395 3063
rect 1565 3037 1612 3043
rect 2276 3036 2278 3044
rect 6010 3036 6012 3044
rect 3112 3006 3113 3014
rect 3121 3006 3123 3014
rect 3131 3006 3133 3014
rect 3141 3006 3143 3014
rect 3151 3006 3160 3014
rect 356 2976 358 2984
rect 1834 2976 1836 2984
rect 3578 2976 3580 2984
rect 5188 2976 5190 2984
rect 164 2917 179 2923
rect 205 2923 211 2943
rect 573 2937 595 2943
rect 836 2937 851 2943
rect 1069 2943 1075 2963
rect 2045 2957 2067 2963
rect 2948 2957 2963 2963
rect 6068 2956 6076 2964
rect 1069 2937 1084 2943
rect 1213 2937 1228 2943
rect 1469 2937 1484 2943
rect 1757 2937 1788 2943
rect 1837 2937 1852 2943
rect 2093 2937 2108 2943
rect 2221 2937 2236 2943
rect 2644 2937 2659 2943
rect 3517 2937 3532 2943
rect 3581 2937 3635 2943
rect 3645 2937 3676 2943
rect 3812 2937 3827 2943
rect 3885 2937 3916 2943
rect 205 2917 227 2923
rect 221 2884 227 2917
rect 637 2917 668 2923
rect 980 2917 995 2923
rect 1053 2917 1068 2923
rect 1421 2917 1436 2923
rect 1581 2917 1628 2923
rect 2324 2917 2355 2923
rect 2365 2917 2380 2923
rect 2637 2917 2643 2936
rect 2781 2917 2787 2936
rect 2941 2917 2956 2923
rect 3085 2917 3164 2923
rect 3389 2917 3404 2923
rect 3789 2917 3820 2923
rect 4157 2923 4163 2943
rect 4972 2943 4980 2948
rect 4564 2937 4595 2943
rect 4765 2937 4804 2943
rect 4972 2937 4995 2943
rect 5028 2937 5043 2943
rect 5085 2937 5123 2943
rect 5949 2937 5980 2943
rect 4157 2917 4211 2923
rect 5005 2917 5043 2923
rect 253 2897 275 2903
rect 429 2897 451 2903
rect 996 2896 1004 2904
rect 2868 2897 2883 2903
rect 3741 2897 3763 2903
rect 5037 2897 5043 2917
rect 5220 2917 5235 2923
rect 5357 2917 5379 2923
rect 5469 2917 5491 2923
rect 5524 2917 5532 2923
rect 5565 2917 5603 2923
rect 5565 2897 5571 2917
rect 5988 2917 6003 2923
rect 252 2884 260 2888
rect 4100 2876 4104 2884
rect 5869 2877 5923 2883
rect 1581 2857 1628 2863
rect 2276 2836 2278 2844
rect 3082 2836 3084 2844
rect 6180 2836 6182 2844
rect 1576 2806 1577 2814
rect 1585 2806 1587 2814
rect 1595 2806 1597 2814
rect 1605 2806 1607 2814
rect 1615 2806 1624 2814
rect 4664 2806 4665 2814
rect 4673 2806 4675 2814
rect 4683 2806 4685 2814
rect 4693 2806 4695 2814
rect 4703 2806 4712 2814
rect 2020 2776 2022 2784
rect 2148 2776 2150 2784
rect 2580 2776 2582 2784
rect 2954 2776 2956 2784
rect 3412 2776 3414 2784
rect 3578 2776 3580 2784
rect 3658 2776 3660 2784
rect 3732 2776 3734 2784
rect 5754 2776 5756 2784
rect 6212 2776 6214 2784
rect 218 2756 220 2764
rect 3956 2756 3960 2764
rect 1156 2736 1158 2744
rect 1828 2736 1830 2744
rect 3012 2736 3014 2744
rect 4042 2736 4044 2744
rect 5588 2736 5590 2744
rect 964 2717 979 2723
rect 1604 2717 1619 2723
rect 1853 2717 1875 2723
rect 3085 2717 3100 2723
rect 317 2697 332 2703
rect 476 2703 484 2708
rect 476 2697 499 2703
rect 493 2684 499 2697
rect 972 2703 980 2708
rect 972 2697 995 2703
rect 1140 2697 1155 2703
rect 1556 2697 1612 2703
rect 1796 2697 1827 2703
rect 2004 2697 2012 2703
rect 2093 2697 2124 2703
rect 2365 2697 2387 2703
rect 157 2677 172 2683
rect 589 2677 627 2683
rect 1549 2677 1619 2683
rect 1972 2677 2003 2683
rect 2173 2677 2195 2683
rect 2285 2677 2307 2683
rect 2509 2677 2515 2716
rect 2541 2697 2556 2703
rect 2541 2684 2547 2697
rect 2669 2697 2684 2703
rect 3117 2697 3148 2703
rect 3117 2684 3123 2697
rect 3284 2697 3299 2703
rect 3309 2697 3324 2703
rect 109 2657 140 2663
rect 2876 2663 2884 2666
rect 1501 2657 1532 2663
rect 1725 2657 1747 2663
rect 2429 2657 2451 2663
rect 2876 2657 2899 2663
rect 3293 2657 3299 2697
rect 4020 2697 4035 2703
rect 4253 2697 4268 2703
rect 4845 2697 4883 2703
rect 5165 2697 5203 2703
rect 5517 2697 5539 2703
rect 5613 2703 5619 2723
rect 5572 2697 5587 2703
rect 5613 2697 5651 2703
rect 5661 2697 5715 2703
rect 5876 2697 5891 2703
rect 5940 2697 5955 2703
rect 5556 2677 5571 2683
rect 5837 2677 5852 2683
rect 6141 2677 6147 2736
rect 6061 2657 6076 2663
rect 2212 2636 2214 2644
rect 4180 2636 4184 2644
rect 3112 2606 3113 2614
rect 3121 2606 3123 2614
rect 3131 2606 3133 2614
rect 3141 2606 3143 2614
rect 3151 2606 3160 2614
rect 3752 2576 3756 2584
rect 5482 2576 5484 2584
rect 1100 2557 1116 2563
rect 1100 2554 1108 2557
rect 1245 2557 1283 2563
rect 1581 2557 1651 2563
rect 1933 2557 1955 2563
rect 4381 2557 4403 2563
rect 4605 2557 4652 2563
rect 173 2537 220 2543
rect 237 2537 275 2543
rect 813 2537 867 2543
rect 1133 2537 1148 2543
rect 1757 2537 1772 2543
rect 2445 2537 2460 2543
rect 2637 2537 2652 2543
rect 2996 2537 3027 2543
rect 3316 2537 3331 2543
rect 196 2517 211 2523
rect 524 2517 540 2523
rect 524 2514 532 2517
rect 557 2517 572 2523
rect 701 2517 716 2523
rect 1444 2497 1459 2503
rect 1501 2483 1507 2523
rect 1684 2517 1692 2523
rect 1773 2517 1788 2523
rect 2052 2517 2067 2523
rect 2685 2517 2700 2523
rect 3076 2517 3091 2523
rect 3325 2517 3331 2537
rect 3693 2523 3699 2543
rect 4052 2537 4067 2543
rect 4317 2537 4332 2543
rect 5421 2543 5427 2563
rect 5421 2537 5452 2543
rect 5732 2537 5747 2543
rect 3661 2517 3699 2523
rect 3837 2517 3852 2523
rect 4020 2517 4035 2523
rect 4068 2517 4083 2523
rect 4132 2517 4147 2523
rect 4493 2517 4524 2523
rect 4557 2517 4595 2523
rect 4644 2517 4691 2523
rect 5277 2517 5315 2523
rect 5357 2517 5379 2523
rect 6036 2517 6051 2523
rect 4084 2496 4092 2504
rect 4148 2496 4156 2504
rect 1501 2477 1516 2483
rect 2020 2477 2035 2483
rect 2394 2476 2396 2484
rect 3092 2476 3094 2484
rect 5764 2476 5766 2484
rect 6052 2476 6054 2484
rect 1348 2456 1350 2464
rect 2826 2456 2828 2464
rect 1576 2406 1577 2414
rect 1585 2406 1587 2414
rect 1595 2406 1597 2414
rect 1605 2406 1607 2414
rect 1615 2406 1624 2414
rect 4664 2406 4665 2414
rect 4673 2406 4675 2414
rect 4683 2406 4685 2414
rect 4693 2406 4695 2414
rect 4703 2406 4712 2414
rect 1370 2376 1372 2384
rect 1428 2376 1430 2384
rect 2842 2376 2844 2384
rect 2986 2376 2988 2384
rect 3572 2376 3574 2384
rect 4324 2376 4326 2384
rect 1306 2356 1308 2364
rect 1229 2337 1244 2343
rect 1501 2343 1507 2363
rect 2634 2356 2636 2364
rect 1501 2337 1516 2343
rect 3818 2336 3820 2344
rect 4164 2336 4166 2344
rect 4388 2336 4390 2344
rect 4477 2337 4524 2343
rect 1796 2317 1811 2323
rect 2180 2316 2188 2324
rect 2589 2317 2611 2323
rect 2770 2316 2780 2324
rect 461 2297 476 2303
rect 564 2297 595 2303
rect 605 2297 636 2303
rect 1309 2297 1324 2303
rect 1373 2297 1388 2303
rect 1396 2297 1427 2303
rect 1773 2297 1788 2303
rect 2637 2297 2675 2303
rect 2845 2297 2876 2303
rect 3437 2297 3459 2303
rect 3789 2303 3795 2323
rect 4477 2317 4483 2337
rect 5197 2337 5212 2343
rect 6260 2336 6262 2344
rect 5244 2332 5252 2336
rect 3757 2297 3795 2303
rect 4269 2297 4307 2303
rect 45 2277 60 2283
rect 365 2277 403 2283
rect 477 2277 499 2283
rect 781 2277 796 2283
rect 628 2257 652 2263
rect 781 2257 787 2277
rect 1396 2277 1411 2283
rect 1828 2277 1843 2283
rect 2701 2277 2716 2283
rect 3380 2277 3395 2283
rect 3860 2277 3875 2283
rect 4301 2277 4307 2297
rect 4932 2297 4947 2303
rect 5085 2297 5116 2303
rect 5652 2297 5667 2303
rect 5757 2303 5763 2323
rect 5725 2297 5763 2303
rect 5789 2297 5820 2303
rect 5981 2303 5987 2323
rect 5981 2297 6019 2303
rect 5004 2277 5028 2283
rect 5981 2277 5996 2283
rect 900 2257 915 2263
rect 1860 2257 1875 2263
rect 708 2236 710 2244
rect 1578 2236 1580 2244
rect 5236 2236 5238 2244
rect 5860 2236 5864 2244
rect 3112 2206 3113 2214
rect 3121 2206 3123 2214
rect 3131 2206 3133 2214
rect 3141 2206 3143 2214
rect 3151 2206 3160 2214
rect 1092 2176 1094 2184
rect 3060 2176 3062 2184
rect 6020 2176 6024 2184
rect 1444 2156 1452 2164
rect 1716 2157 1731 2163
rect 3245 2157 3268 2163
rect 285 2137 307 2143
rect 413 2137 428 2143
rect 237 2117 268 2123
rect 276 2117 291 2123
rect 308 2117 323 2123
rect 749 2117 787 2123
rect 324 2096 332 2104
rect 724 2096 732 2104
rect 749 2097 755 2117
rect 1021 2117 1027 2156
rect 3260 2154 3268 2157
rect 1325 2137 1356 2143
rect 1588 2137 1651 2143
rect 2461 2137 2492 2143
rect 1229 2117 1283 2123
rect 1348 2117 1363 2123
rect 2244 2117 2259 2123
rect 2445 2117 2460 2123
rect 2621 2117 2652 2123
rect 2797 2123 2803 2143
rect 3124 2137 3171 2143
rect 3533 2143 3539 2163
rect 3828 2156 3836 2164
rect 5644 2157 5676 2163
rect 5644 2148 5652 2157
rect 3524 2137 3539 2143
rect 3549 2137 3571 2143
rect 3741 2137 3779 2143
rect 4212 2137 4227 2143
rect 4541 2137 4579 2143
rect 4596 2137 4611 2143
rect 4941 2137 4979 2143
rect 2797 2117 2812 2123
rect 2925 2117 2940 2123
rect 3172 2117 3180 2123
rect 3517 2117 3532 2123
rect 3661 2117 3692 2123
rect 3812 2117 3827 2123
rect 980 2097 995 2103
rect 1005 2083 1011 2103
rect 3821 2097 3827 2117
rect 4781 2117 4819 2123
rect 3906 2096 3916 2104
rect 4493 2097 4515 2103
rect 4781 2097 4787 2117
rect 4884 2117 4899 2123
rect 5476 2117 5507 2123
rect 5869 2123 5875 2143
rect 5860 2117 5875 2123
rect 5981 2123 5987 2143
rect 5981 2117 6012 2123
rect 5101 2097 5139 2103
rect 973 2077 1011 2083
rect 973 2057 979 2077
rect 1485 2077 1539 2083
rect 836 2036 838 2044
rect 1576 2006 1577 2014
rect 1585 2006 1587 2014
rect 1595 2006 1597 2014
rect 1605 2006 1607 2014
rect 1615 2006 1624 2014
rect 4664 2006 4665 2014
rect 4673 2006 4675 2014
rect 4683 2006 4685 2014
rect 4693 2006 4695 2014
rect 4703 2006 4712 2014
rect 1156 1976 1158 1984
rect 2052 1976 2054 1984
rect 3076 1976 3078 1984
rect 3786 1976 3788 1984
rect 3844 1976 3846 1984
rect 4916 1976 4918 1984
rect 4986 1976 4988 1984
rect 5044 1976 5046 1984
rect 6058 1976 6060 1984
rect 5172 1956 5174 1964
rect 1284 1936 1286 1944
rect 3709 1937 3724 1943
rect 4260 1936 4262 1944
rect 5242 1936 5244 1944
rect 5508 1936 5514 1944
rect 6116 1936 6118 1944
rect 6212 1937 6227 1943
rect 4300 1932 4308 1936
rect 292 1916 302 1924
rect 1965 1917 1980 1923
rect 3229 1917 3267 1923
rect 4196 1916 4204 1924
rect 4285 1917 4307 1923
rect 604 1904 612 1908
rect 317 1897 348 1903
rect 1005 1897 1020 1903
rect 1140 1897 1155 1903
rect 1332 1897 1347 1903
rect 1389 1884 1395 1903
rect 1581 1897 1644 1903
rect 237 1877 275 1883
rect 1021 1877 1043 1883
rect 1620 1877 1651 1883
rect 1693 1864 1699 1903
rect 1853 1897 1875 1903
rect 1908 1897 1939 1903
rect 2164 1897 2179 1903
rect 1901 1877 1916 1883
rect 1901 1857 1907 1877
rect 2141 1877 2156 1883
rect 1988 1857 2003 1863
rect 2189 1863 2195 1903
rect 3101 1897 3180 1903
rect 3309 1897 3363 1903
rect 3373 1897 3388 1903
rect 3789 1897 3804 1903
rect 3876 1897 3891 1903
rect 3901 1897 3932 1903
rect 4052 1897 4067 1903
rect 4077 1897 4108 1903
rect 4692 1897 4723 1903
rect 4820 1897 4851 1903
rect 4900 1897 4908 1903
rect 5140 1897 5171 1903
rect 5252 1897 5299 1903
rect 5556 1897 5587 1903
rect 5965 1897 5980 1903
rect 6068 1897 6115 1903
rect 2269 1877 2284 1883
rect 2445 1877 2499 1883
rect 2900 1877 2931 1883
rect 2964 1877 2979 1883
rect 3156 1877 3187 1883
rect 3444 1877 3459 1883
rect 3485 1877 3523 1883
rect 2189 1857 2204 1863
rect 2820 1857 2835 1863
rect 3412 1857 3427 1863
rect 3453 1857 3459 1877
rect 4772 1877 4803 1883
rect 4884 1877 4899 1883
rect 5268 1877 5283 1883
rect 5644 1877 5676 1883
rect 573 1837 588 1843
rect 3594 1836 3596 1844
rect 3112 1806 3113 1814
rect 3121 1806 3123 1814
rect 3131 1806 3133 1814
rect 3141 1806 3143 1814
rect 3151 1806 3160 1814
rect 218 1776 220 1784
rect 628 1776 630 1784
rect 2404 1776 2406 1784
rect 4890 1776 4892 1784
rect 5610 1776 5612 1784
rect 765 1757 780 1763
rect 836 1757 851 1763
rect 428 1743 436 1748
rect 1741 1744 1747 1763
rect 2340 1757 2355 1763
rect 428 1737 451 1743
rect 541 1737 579 1743
rect 596 1737 611 1743
rect 461 1717 499 1723
rect 605 1717 611 1737
rect 653 1737 684 1743
rect 1380 1737 1395 1743
rect 1645 1737 1676 1743
rect 1869 1737 1900 1743
rect 2260 1737 2275 1743
rect 2413 1737 2428 1743
rect 1244 1724 1252 1728
rect 772 1717 835 1723
rect 884 1717 915 1723
rect 1485 1723 1491 1736
rect 2413 1724 2419 1737
rect 2468 1737 2499 1743
rect 1485 1717 1508 1723
rect 1500 1712 1508 1717
rect 61 1697 83 1703
rect 500 1696 508 1704
rect 1517 1684 1523 1723
rect 1549 1717 1596 1723
rect 1885 1717 1900 1723
rect 2141 1717 2179 1723
rect 2228 1717 2243 1723
rect 2637 1717 2643 1756
rect 2669 1724 2675 1763
rect 2781 1757 2808 1763
rect 3485 1737 3500 1743
rect 3773 1737 3811 1743
rect 3236 1717 3251 1723
rect 3549 1717 3564 1723
rect 3661 1717 3692 1723
rect 3773 1717 3779 1737
rect 5140 1737 5148 1743
rect 5741 1737 5763 1743
rect 4333 1717 4371 1723
rect 4749 1717 4787 1723
rect 1466 1676 1468 1684
rect 1789 1683 1795 1703
rect 3485 1697 3507 1703
rect 3677 1697 3715 1703
rect 4724 1696 4732 1704
rect 4749 1697 4755 1717
rect 4845 1717 4860 1723
rect 5076 1717 5091 1723
rect 5140 1717 5171 1723
rect 5181 1717 5219 1723
rect 5245 1717 5260 1723
rect 5213 1697 5219 1717
rect 5501 1717 5539 1723
rect 5565 1717 5580 1723
rect 5236 1696 5244 1704
rect 5533 1697 5539 1717
rect 5764 1717 5779 1723
rect 1773 1677 1795 1683
rect 3882 1656 3884 1664
rect 4637 1657 4652 1663
rect 5844 1656 5846 1664
rect 1268 1636 1270 1644
rect 1572 1637 1596 1643
rect 2292 1636 2294 1644
rect 2708 1636 2710 1644
rect 3588 1636 3590 1644
rect 3764 1636 3766 1644
rect 4420 1636 4422 1644
rect 4842 1636 4844 1644
rect 1576 1606 1577 1614
rect 1585 1606 1587 1614
rect 1595 1606 1597 1614
rect 1605 1606 1607 1614
rect 1615 1606 1624 1614
rect 4664 1606 4665 1614
rect 4673 1606 4675 1614
rect 4683 1606 4685 1614
rect 4693 1606 4695 1614
rect 4703 1606 4712 1614
rect 436 1576 438 1584
rect 1396 1576 1398 1584
rect 1700 1576 1702 1584
rect 2266 1576 2268 1584
rect 5812 1576 5814 1584
rect 100 1537 115 1543
rect 1117 1537 1132 1543
rect 2493 1543 2499 1563
rect 2493 1537 2508 1543
rect 4250 1536 4252 1544
rect 4676 1537 4732 1543
rect 6010 1536 6012 1544
rect 4380 1532 4388 1536
rect 36 1516 44 1524
rect 45 1497 83 1503
rect 461 1503 467 1523
rect 557 1517 595 1523
rect 868 1516 876 1524
rect 461 1497 483 1503
rect 340 1477 371 1483
rect 477 1483 483 1497
rect 717 1497 732 1503
rect 477 1477 499 1483
rect 717 1457 723 1497
rect 813 1497 844 1503
rect 1469 1483 1475 1503
rect 1661 1497 1676 1503
rect 1444 1477 1459 1483
rect 1469 1477 1484 1483
rect 1533 1477 1548 1483
rect 1661 1477 1667 1497
rect 1725 1503 1731 1523
rect 1917 1517 1939 1523
rect 2612 1517 2627 1523
rect 1725 1497 1747 1503
rect 1741 1484 1747 1497
rect 2093 1497 2156 1503
rect 2404 1497 2412 1503
rect 2644 1497 2668 1503
rect 2861 1497 2876 1503
rect 2909 1497 2940 1503
rect 3124 1497 3139 1503
rect 3620 1497 3651 1503
rect 3965 1503 3971 1523
rect 4148 1516 4156 1524
rect 4205 1517 4227 1523
rect 4333 1517 4371 1523
rect 4669 1517 4684 1523
rect 3933 1497 3971 1503
rect 4292 1497 4307 1503
rect 4781 1503 4787 1523
rect 5300 1516 5308 1524
rect 4749 1497 4787 1503
rect 5332 1497 5363 1503
rect 5556 1497 5587 1503
rect 5709 1497 5724 1503
rect 2148 1477 2163 1483
rect 2644 1477 2675 1483
rect 2868 1477 2883 1483
rect 3613 1477 3628 1483
rect 3956 1477 3971 1483
rect 5389 1477 5420 1483
rect 5709 1483 5715 1497
rect 5732 1497 5740 1503
rect 5844 1497 5875 1503
rect 6036 1497 6067 1503
rect 5693 1477 5715 1483
rect 5484 1472 5492 1476
rect 1421 1457 1443 1463
rect 1549 1457 1564 1463
rect 3044 1456 3052 1464
rect 3468 1463 3476 1466
rect 3468 1457 3491 1463
rect 1288 1436 1292 1444
rect 1572 1437 1619 1443
rect 1908 1436 1910 1444
rect 3092 1437 3100 1443
rect 3112 1406 3113 1414
rect 3121 1406 3123 1414
rect 3131 1406 3133 1414
rect 3141 1406 3143 1414
rect 3151 1406 3160 1414
rect 1130 1376 1132 1384
rect 2205 1377 2243 1383
rect 2237 1364 2243 1377
rect 3332 1376 3336 1384
rect 4605 1377 4620 1383
rect 420 1357 435 1363
rect 1620 1357 1667 1363
rect 3037 1357 3052 1363
rect 4828 1344 4836 1348
rect 52 1337 60 1343
rect 141 1337 188 1343
rect 381 1337 412 1343
rect 797 1337 812 1343
rect 1540 1337 1555 1343
rect 1597 1337 1644 1343
rect 2116 1337 2131 1343
rect 2381 1337 2396 1343
rect 324 1317 371 1323
rect 660 1317 675 1323
rect 733 1317 771 1323
rect 797 1317 835 1323
rect 797 1297 803 1317
rect 1092 1317 1123 1323
rect 1197 1317 1212 1323
rect 1117 1297 1123 1317
rect 1332 1317 1347 1323
rect 1556 1317 1571 1323
rect 1764 1317 1788 1323
rect 2413 1323 2419 1343
rect 2509 1337 2524 1343
rect 3213 1337 3244 1343
rect 3661 1337 3683 1343
rect 3949 1337 3971 1343
rect 5028 1337 5059 1343
rect 5405 1337 5420 1343
rect 5428 1337 5443 1343
rect 2404 1317 2419 1323
rect 2621 1317 2636 1323
rect 2804 1317 2812 1323
rect 2893 1317 2947 1323
rect 3684 1317 3699 1323
rect 3972 1317 3987 1323
rect 4036 1317 4051 1323
rect 4356 1317 4371 1323
rect 4532 1317 4547 1323
rect 4733 1317 4764 1323
rect 5140 1317 5155 1323
rect 5284 1317 5299 1323
rect 5469 1317 5507 1323
rect 1508 1296 1516 1304
rect 3700 1296 3708 1304
rect 3988 1296 3996 1304
rect 4386 1296 4396 1304
rect 4884 1296 4892 1304
rect 5501 1297 5507 1317
rect 4845 1277 4868 1283
rect 6116 1276 6122 1284
rect 1754 1236 1756 1244
rect 2436 1236 2438 1244
rect 1576 1206 1577 1214
rect 1585 1206 1587 1214
rect 1595 1206 1597 1214
rect 1605 1206 1607 1214
rect 1615 1206 1624 1214
rect 4664 1206 4665 1214
rect 4673 1206 4675 1214
rect 4683 1206 4685 1214
rect 4693 1206 4695 1214
rect 4703 1206 4712 1214
rect 1876 1176 1878 1184
rect 4970 1176 4972 1184
rect 5028 1176 5030 1184
rect 5732 1176 5734 1184
rect 5866 1176 5868 1184
rect 6228 1176 6230 1184
rect 493 1137 508 1143
rect 676 1137 684 1143
rect 973 1137 988 1143
rect 3004 1137 3027 1143
rect 4109 1137 4124 1143
rect 4324 1137 4339 1143
rect 109 1097 124 1103
rect 157 1097 172 1103
rect 301 1097 316 1103
rect 349 1097 403 1103
rect 893 1103 899 1123
rect 948 1117 963 1123
rect 996 1117 1011 1123
rect 1044 1117 1059 1123
rect 836 1097 867 1103
rect 893 1097 908 1103
rect 1133 1103 1139 1136
rect 2396 1124 2404 1128
rect 1325 1117 1340 1123
rect 1492 1117 1507 1123
rect 2429 1117 2444 1123
rect 2877 1117 2899 1123
rect 1133 1097 1155 1103
rect 436 1077 451 1083
rect 1149 1077 1155 1097
rect 1421 1097 1436 1103
rect 1837 1097 1875 1103
rect 1892 1097 1900 1103
rect 2884 1097 2899 1103
rect 3124 1097 3164 1103
rect 3421 1103 3427 1123
rect 3389 1097 3427 1103
rect 3508 1097 3523 1103
rect 3828 1097 3843 1103
rect 4141 1097 4163 1103
rect 4372 1097 4387 1103
rect 1556 1077 1571 1083
rect 2260 1077 2275 1083
rect 2573 1077 2611 1083
rect 2836 1077 2844 1083
rect 4349 1083 4355 1096
rect 4349 1077 4371 1083
rect 253 1057 268 1063
rect 1693 1057 1708 1063
rect 2781 1057 2819 1063
rect 3501 1057 3516 1063
rect 4365 1057 4371 1077
rect 4397 1064 4403 1103
rect 4765 1097 4819 1103
rect 4852 1097 4867 1103
rect 4973 1097 4988 1103
rect 5037 1097 5075 1103
rect 5085 1097 5100 1103
rect 5421 1103 5427 1123
rect 5652 1117 5667 1123
rect 5380 1097 5411 1103
rect 5421 1097 5436 1103
rect 5444 1097 5459 1103
rect 5677 1097 5708 1103
rect 5869 1097 5884 1103
rect 6100 1097 6115 1103
rect 4669 1077 4684 1083
rect 4909 1077 4924 1083
rect 5332 1077 5363 1083
rect 5581 1077 5596 1083
rect 5917 1077 5955 1083
rect 6196 1077 6211 1083
rect 5197 1057 5235 1063
rect 5972 1057 5996 1063
rect 1018 1036 1020 1044
rect 1924 1036 1926 1044
rect 3117 1037 3164 1043
rect 4708 1037 4739 1043
rect 6052 1036 6054 1044
rect 3112 1006 3113 1014
rect 3121 1006 3123 1014
rect 3131 1006 3133 1014
rect 3141 1006 3143 1014
rect 3151 1006 3160 1014
rect 84 976 86 984
rect 170 976 172 984
rect 1178 976 1180 984
rect 3028 977 3043 983
rect 4132 976 4134 984
rect 5540 976 5542 984
rect 132 956 140 964
rect 404 957 419 963
rect 500 957 515 963
rect 100 937 115 943
rect 237 937 252 943
rect 285 937 300 943
rect 685 943 691 963
rect 932 957 947 963
rect 1604 957 1644 963
rect 685 937 700 943
rect 916 937 931 943
rect 397 917 412 923
rect 708 917 723 923
rect 925 917 931 937
rect 1028 937 1043 943
rect 1133 937 1164 943
rect 2045 943 2051 963
rect 2356 957 2371 963
rect 2541 957 2556 963
rect 4877 957 4892 963
rect 4909 957 4924 963
rect 5636 956 5644 964
rect 5917 957 5932 963
rect 1844 937 1875 943
rect 2045 937 2060 943
rect 2148 937 2163 943
rect 2429 937 2460 943
rect 2596 937 2627 943
rect 4589 937 4604 943
rect 4836 937 4851 943
rect 5053 937 5091 943
rect 1620 917 1660 923
rect 1821 917 1836 923
rect 1997 917 2019 923
rect 2189 917 2220 923
rect 2276 917 2307 923
rect 2477 917 2492 923
rect 2548 917 2563 923
rect 2829 917 2844 923
rect 2909 917 2947 923
rect 45 897 60 903
rect 141 897 156 903
rect 244 897 259 903
rect 429 897 451 903
rect 628 897 643 903
rect 1069 897 1091 903
rect 1149 897 1164 903
rect 1300 897 1315 903
rect 1508 896 1516 904
rect 1917 897 1932 903
rect 2269 897 2284 903
rect 2941 897 2947 917
rect 3549 917 3564 923
rect 4925 917 4963 923
rect 5037 917 5052 923
rect 5236 917 5251 923
rect 5341 923 5347 943
rect 5444 937 5459 943
rect 5613 937 5651 943
rect 5972 937 5980 943
rect 5284 917 5315 923
rect 5341 917 5356 923
rect 5549 917 5564 923
rect 5549 897 5555 917
rect 5988 917 5996 923
rect 6269 917 6307 923
rect 44 884 52 888
rect 6301 884 6307 917
rect 628 877 659 883
rect 1277 877 1292 883
rect 1277 857 1283 877
rect 1325 877 1340 883
rect 3012 877 3043 883
rect 5252 876 5254 884
rect 5421 877 5436 883
rect 1380 856 1382 864
rect 2026 856 2028 864
rect 724 836 726 844
rect 1684 836 1686 844
rect 1818 836 1820 844
rect 2244 836 2246 844
rect 4570 836 4572 844
rect 1576 806 1577 814
rect 1585 806 1587 814
rect 1595 806 1597 814
rect 1605 806 1607 814
rect 1615 806 1624 814
rect 4664 806 4665 814
rect 4673 806 4675 814
rect 4683 806 4685 814
rect 4693 806 4695 814
rect 4703 806 4712 814
rect 186 776 188 784
rect 506 776 508 784
rect 2842 776 2844 784
rect 4004 776 4006 784
rect 4858 776 4860 784
rect 5364 776 5366 784
rect 6100 776 6102 784
rect 3620 756 3622 764
rect 4653 757 4707 763
rect 45 737 60 743
rect 973 737 1012 743
rect 621 717 636 723
rect 77 697 92 703
rect 157 697 179 703
rect 237 697 259 703
rect 333 697 348 703
rect 365 697 387 703
rect 973 697 979 737
rect 1434 736 1436 744
rect 1492 736 1494 744
rect 1629 737 1644 743
rect 3901 737 3924 743
rect 1517 717 1555 723
rect 1565 717 1635 723
rect 1037 697 1052 703
rect 1261 697 1292 703
rect 1341 697 1372 703
rect 1709 703 1715 723
rect 1709 697 1747 703
rect 2045 703 2051 723
rect 2013 697 2051 703
rect 2276 697 2307 703
rect 2477 703 2483 723
rect 3117 717 3132 723
rect 2404 697 2435 703
rect 2445 697 2483 703
rect 2532 697 2572 703
rect 2676 697 2691 703
rect 2749 697 2764 703
rect 2868 697 2899 703
rect 2996 697 3011 703
rect 420 677 444 683
rect 628 677 643 683
rect 952 676 956 684
rect 1213 677 1244 683
rect 1293 677 1299 696
rect 1389 677 1420 683
rect 1453 677 1475 683
rect 1453 664 1459 677
rect 1572 677 1612 683
rect 2381 677 2419 683
rect 2525 677 2531 696
rect 2564 677 2579 683
rect 3373 677 3404 683
rect 3485 683 3491 736
rect 4653 723 4659 757
rect 4749 743 4755 763
rect 4724 737 4755 743
rect 5885 737 5939 743
rect 4612 717 4627 723
rect 4637 717 4659 723
rect 5069 717 5091 723
rect 3604 697 3619 703
rect 3901 697 3916 703
rect 4189 697 4204 703
rect 4365 692 4371 716
rect 4388 697 4403 703
rect 4436 697 4451 703
rect 3453 677 3491 683
rect 3501 677 3539 683
rect 3709 677 3724 683
rect 3796 677 3827 683
rect 3965 677 3980 683
rect 4196 677 4211 683
rect 4244 677 4252 683
rect 4365 677 4380 683
rect 4445 677 4451 697
rect 4532 697 4547 703
rect 4644 697 4684 703
rect 4932 697 4963 703
rect 4973 697 5004 703
rect 5469 684 5475 703
rect 5636 697 5651 703
rect 5773 697 5788 703
rect 5885 697 5891 737
rect 5933 697 5948 703
rect 6109 697 6147 703
rect 6164 697 6195 703
rect 4644 677 4668 683
rect 5284 677 5292 683
rect 5556 677 5564 683
rect 5629 677 5644 683
rect 132 657 147 663
rect 285 657 300 663
rect 4500 657 4515 663
rect 554 636 556 644
rect 2794 636 2796 644
rect 3252 636 3254 644
rect 3300 636 3302 644
rect 3562 636 3564 644
rect 4228 636 4230 644
rect 4468 636 4470 644
rect 4637 637 4684 643
rect 3112 606 3113 614
rect 3121 606 3123 614
rect 3131 606 3133 614
rect 3141 606 3143 614
rect 3151 606 3160 614
rect 1130 576 1132 584
rect 5048 576 5052 584
rect 333 557 348 563
rect 1172 557 1187 563
rect 461 537 492 543
rect 1053 537 1107 543
rect 1396 537 1411 543
rect 1533 543 1539 563
rect 1645 557 1667 563
rect 3572 556 3580 564
rect 3629 557 3644 563
rect 1524 537 1539 543
rect 1780 537 1795 543
rect 2340 537 2348 543
rect 2365 537 2380 543
rect 2500 537 2515 543
rect 2701 537 2739 543
rect 2877 537 2908 543
rect 2941 537 2956 543
rect 3101 537 3164 543
rect 3325 537 3340 543
rect 397 517 451 523
rect 717 517 764 523
rect 868 517 883 523
rect 1181 517 1235 523
rect 1261 517 1299 523
rect 797 497 835 503
rect 1261 497 1267 517
rect 1412 517 1427 523
rect 1565 517 1580 523
rect 2141 517 2179 523
rect 1940 496 1948 504
rect 2173 497 2179 517
rect 2557 517 2595 523
rect 2605 517 2620 523
rect 2429 497 2451 503
rect 2557 497 2563 517
rect 3012 517 3036 523
rect 3293 517 3315 523
rect 3581 517 3596 523
rect 3044 496 3052 504
rect 3156 497 3180 503
rect 3229 497 3251 503
rect 906 476 908 484
rect 3469 483 3475 503
rect 3581 497 3587 517
rect 3629 517 3635 557
rect 4148 557 4163 563
rect 4573 557 4588 563
rect 5197 557 5228 563
rect 5908 557 5923 563
rect 3677 543 3683 556
rect 3677 537 3699 543
rect 4068 537 4099 543
rect 4660 537 4723 543
rect 4884 537 4899 543
rect 4932 537 4963 543
rect 5220 537 5251 543
rect 5492 537 5507 543
rect 5668 537 5676 543
rect 4397 517 4412 523
rect 5172 517 5203 523
rect 5220 517 5235 523
rect 5245 517 5283 523
rect 5405 517 5443 523
rect 5533 517 5548 523
rect 3885 497 3907 503
rect 4765 497 4780 503
rect 5277 497 5283 517
rect 6084 517 6099 523
rect 3469 477 3516 483
rect 6004 476 6006 484
rect 1565 457 1612 463
rect 1370 436 1372 444
rect 1428 436 1430 444
rect 1738 436 1740 444
rect 1892 436 1894 444
rect 2314 436 2316 444
rect 2532 436 2534 444
rect 2756 436 2758 444
rect 2980 436 2982 444
rect 3620 436 3622 444
rect 3716 436 3718 444
rect 3796 436 3798 444
rect 4858 436 4860 444
rect 5338 436 5340 444
rect 1576 406 1577 414
rect 1585 406 1587 414
rect 1595 406 1597 414
rect 1605 406 1607 414
rect 1615 406 1624 414
rect 4664 406 4665 414
rect 4673 406 4675 414
rect 4683 406 4685 414
rect 4693 406 4695 414
rect 4703 406 4712 414
rect 5194 376 5196 384
rect 2468 356 2470 364
rect 1236 337 1251 343
rect 1652 336 1654 344
rect 2820 337 2851 343
rect 3549 343 3555 363
rect 4090 356 4092 364
rect 4276 356 4278 364
rect 3540 337 3555 343
rect 3620 336 3622 344
rect 6141 337 6195 343
rect 1101 303 1107 323
rect 1892 316 1900 324
rect 4365 317 4403 323
rect 4692 317 4739 323
rect 6084 316 6092 324
rect 1101 297 1139 303
rect 1508 297 1539 303
rect 1572 297 1651 303
rect 1709 297 1724 303
rect 2004 297 2019 303
rect 2093 297 2115 303
rect 1172 277 1187 283
rect 1181 257 1187 277
rect 2276 277 2291 283
rect 2436 277 2451 283
rect 2701 277 2732 283
rect 1197 257 1235 263
rect 1565 257 1612 263
rect 2036 257 2051 263
rect 2628 257 2643 263
rect 2813 244 2819 303
rect 3085 297 3219 303
rect 3428 297 3443 303
rect 3476 297 3491 303
rect 3501 297 3516 303
rect 3741 297 3756 303
rect 4420 297 4451 303
rect 5268 297 5283 303
rect 5588 297 5596 303
rect 5652 297 5667 303
rect 2909 277 2924 283
rect 3101 277 3132 283
rect 3316 277 3331 283
rect 3469 277 3484 283
rect 3972 277 3987 283
rect 4653 277 4684 283
rect 4957 277 4972 283
rect 5572 277 5603 283
rect 5741 283 5747 303
rect 6093 297 6108 303
rect 5732 277 5747 283
rect 5757 277 5788 283
rect 3325 257 3340 263
rect 4564 257 4579 263
rect 5245 257 5260 263
rect 5837 257 5852 263
rect 1092 236 1094 244
rect 1976 236 1980 244
rect 2948 236 2952 244
rect 3668 237 3683 243
rect 3944 236 3948 244
rect 4356 236 4358 244
rect 4776 236 4780 244
rect 4996 236 4998 244
rect 5492 237 5507 243
rect 3112 206 3113 214
rect 3121 206 3123 214
rect 3131 206 3133 214
rect 3141 206 3143 214
rect 3151 206 3160 214
rect 3700 176 3702 184
rect 6004 176 6006 184
rect 1437 157 1468 163
rect 1716 157 1731 163
rect 1741 157 1756 163
rect 2104 156 2108 164
rect 2445 157 2460 163
rect 1284 137 1299 143
rect 1620 137 1644 143
rect 2508 143 2516 144
rect 2500 137 2516 143
rect 2637 143 2643 163
rect 3117 157 3196 163
rect 3252 157 3267 163
rect 3416 157 3443 163
rect 4477 144 4483 163
rect 4804 157 4819 163
rect 4829 157 4860 163
rect 2637 137 2652 143
rect 764 117 803 123
rect 764 116 772 117
rect 916 117 947 123
rect 1149 117 1187 123
rect 1261 117 1292 123
rect 1181 97 1187 117
rect 1597 117 1660 123
rect 1757 117 1779 123
rect 1997 117 2019 123
rect 2685 123 2691 143
rect 3124 137 3196 143
rect 3261 137 3276 143
rect 3476 137 3507 143
rect 3517 137 3532 143
rect 3885 137 3916 143
rect 4205 137 4236 143
rect 4269 137 4323 143
rect 4429 137 4444 143
rect 4813 137 4828 143
rect 4957 137 4972 143
rect 5076 137 5091 143
rect 6093 137 6108 143
rect 2589 117 2611 123
rect 2621 117 2659 123
rect 2685 117 2707 123
rect 1965 97 1980 103
rect 2653 97 2659 117
rect 2845 117 2883 123
rect 3069 117 3091 123
rect 3597 117 3619 123
rect 3933 117 3964 123
rect 3997 117 4019 123
rect 4084 117 4099 123
rect 4116 117 4124 123
rect 4173 117 4211 123
rect 4228 117 4243 123
rect 4532 117 4563 123
rect 4628 117 4643 123
rect 4797 117 4812 123
rect 3037 97 3052 103
rect 3709 97 3731 103
rect 3780 97 3795 103
rect 4637 97 4643 117
rect 4877 117 4915 123
rect 4909 97 4915 117
rect 5021 117 5059 123
rect 4932 96 4940 104
rect 5021 97 5027 117
rect 5284 117 5299 123
rect 5293 97 5299 117
rect 5437 97 5452 103
rect 884 76 886 84
rect 1050 76 1052 84
rect 1117 77 1132 83
rect 2026 76 2028 84
rect 3357 77 3411 83
rect 2884 36 2886 44
rect 3460 36 3462 44
rect 1576 6 1577 14
rect 1585 6 1587 14
rect 1595 6 1597 14
rect 1605 6 1607 14
rect 1615 6 1624 14
rect 4664 6 4665 14
rect 4673 6 4675 14
rect 4683 6 4685 14
rect 4693 6 4695 14
rect 4703 6 4712 14
<< m2contact >>
rect 3113 4606 3121 4614
rect 3123 4606 3131 4614
rect 3133 4606 3141 4614
rect 3143 4606 3151 4614
rect 156 4576 164 4584
rect 588 4576 596 4584
rect 748 4576 756 4584
rect 972 4576 980 4584
rect 1164 4576 1172 4584
rect 1388 4576 1396 4584
rect 1724 4576 1732 4584
rect 1900 4576 1908 4584
rect 1948 4576 1956 4584
rect 1964 4576 1972 4584
rect 2012 4576 2020 4584
rect 2092 4576 2100 4584
rect 2284 4576 2292 4584
rect 2444 4576 2452 4584
rect 2636 4576 2644 4584
rect 2796 4576 2804 4584
rect 3020 4576 3028 4584
rect 3068 4576 3076 4584
rect 3692 4576 3700 4584
rect 4060 4576 4068 4584
rect 4444 4576 4452 4584
rect 4828 4576 4836 4584
rect 6236 4576 6244 4584
rect 140 4556 148 4564
rect 604 4556 612 4564
rect 988 4556 996 4564
rect 1148 4556 1156 4564
rect 1372 4556 1380 4564
rect 1804 4556 1812 4564
rect 2428 4556 2436 4564
rect 2732 4556 2740 4564
rect 3036 4556 3044 4564
rect 3052 4556 3060 4564
rect 3676 4556 3684 4564
rect 4092 4556 4100 4564
rect 4428 4556 4436 4564
rect 4700 4556 4708 4564
rect 5788 4556 5796 4564
rect 6060 4556 6068 4564
rect 6092 4556 6100 4564
rect 44 4536 52 4544
rect 108 4536 116 4544
rect 268 4536 276 4544
rect 460 4536 468 4544
rect 668 4536 676 4544
rect 732 4536 740 4544
rect 844 4536 852 4544
rect 1020 4536 1028 4544
rect 1068 4536 1076 4544
rect 1276 4536 1284 4544
rect 1372 4536 1380 4544
rect 1500 4536 1508 4544
rect 1580 4536 1588 4544
rect 1612 4536 1620 4544
rect 1788 4536 1796 4544
rect 1804 4536 1812 4544
rect 2172 4536 2180 4544
rect 2300 4536 2308 4544
rect 2396 4536 2404 4544
rect 2556 4536 2564 4544
rect 2684 4536 2692 4544
rect 2780 4536 2788 4544
rect 2908 4536 2916 4544
rect 3276 4536 3284 4544
rect 3356 4536 3364 4544
rect 3420 4536 3428 4544
rect 3452 4536 3460 4544
rect 3516 4536 3524 4544
rect 3948 4536 3956 4544
rect 4140 4536 4148 4544
rect 4204 4536 4212 4544
rect 4348 4536 4356 4544
rect 4572 4536 4580 4544
rect 4716 4536 4724 4544
rect 4780 4536 4788 4544
rect 4812 4536 4820 4544
rect 4956 4536 4964 4544
rect 5244 4536 5252 4544
rect 5372 4536 5380 4544
rect 5436 4536 5444 4544
rect 5532 4536 5540 4544
rect 5548 4536 5556 4544
rect 5868 4536 5876 4544
rect 5884 4536 5892 4544
rect 5932 4536 5940 4544
rect 5948 4536 5956 4544
rect 5996 4536 6004 4544
rect 6092 4536 6100 4544
rect 6156 4536 6164 4544
rect 6188 4536 6196 4544
rect 6284 4536 6292 4544
rect 252 4516 260 4524
rect 396 4516 404 4524
rect 476 4516 484 4524
rect 668 4516 676 4524
rect 716 4516 724 4524
rect 780 4516 788 4524
rect 860 4516 868 4524
rect 1084 4516 1092 4524
rect 1100 4516 1108 4524
rect 1260 4516 1268 4524
rect 1516 4518 1524 4526
rect 1628 4516 1636 4524
rect 1692 4516 1700 4524
rect 1740 4516 1748 4524
rect 1788 4516 1796 4524
rect 1916 4516 1924 4524
rect 1996 4516 2004 4524
rect 2044 4516 2052 4524
rect 2060 4516 2068 4524
rect 2204 4516 2212 4524
rect 2300 4516 2308 4524
rect 2572 4518 2580 4526
rect 12 4496 20 4504
rect 92 4496 100 4504
rect 620 4496 628 4504
rect 636 4496 644 4504
rect 1020 4496 1028 4504
rect 1052 4496 1060 4504
rect 1116 4496 1124 4504
rect 1644 4496 1652 4504
rect 1676 4496 1684 4504
rect 1740 4496 1748 4504
rect 2316 4496 2324 4504
rect 2668 4516 2676 4524
rect 2364 4496 2372 4504
rect 2716 4496 2724 4504
rect 2764 4516 2772 4524
rect 2892 4518 2900 4526
rect 3100 4516 3108 4524
rect 3260 4516 3268 4524
rect 3372 4516 3380 4524
rect 3532 4516 3540 4524
rect 3804 4516 3812 4524
rect 3964 4516 3972 4524
rect 3420 4496 3428 4504
rect 4140 4496 4148 4504
rect 4204 4516 4212 4524
rect 4332 4516 4340 4524
rect 4540 4516 4548 4524
rect 4636 4516 4644 4524
rect 4732 4516 4740 4524
rect 4940 4516 4948 4524
rect 5020 4516 5028 4524
rect 5260 4518 5268 4526
rect 5324 4516 5332 4524
rect 5356 4516 5364 4524
rect 5420 4516 5428 4524
rect 5580 4516 5588 4524
rect 5612 4516 5620 4524
rect 5692 4516 5700 4524
rect 5740 4516 5748 4524
rect 5916 4516 5924 4524
rect 5932 4516 5940 4524
rect 6012 4516 6020 4524
rect 6060 4516 6068 4524
rect 6108 4516 6116 4524
rect 6172 4516 6180 4524
rect 6204 4516 6212 4524
rect 4780 4496 4788 4504
rect 5100 4496 5108 4504
rect 5116 4496 5124 4504
rect 5324 4496 5332 4504
rect 5388 4496 5396 4504
rect 5420 4496 5428 4504
rect 5452 4496 5460 4504
rect 5500 4496 5508 4504
rect 5580 4496 5588 4504
rect 5596 4496 5604 4504
rect 5708 4496 5716 4504
rect 5788 4496 5796 4504
rect 5836 4496 5844 4504
rect 5884 4496 5892 4504
rect 5980 4496 5988 4504
rect 6044 4496 6052 4504
rect 6236 4496 6244 4504
rect 1036 4476 1044 4484
rect 3164 4476 3172 4484
rect 3676 4476 3684 4484
rect 4860 4476 4868 4484
rect 5628 4476 5636 4484
rect 5660 4476 5668 4484
rect 5676 4476 5684 4484
rect 5756 4476 5764 4484
rect 6012 4476 6020 4484
rect 6300 4476 6308 4484
rect 364 4456 372 4464
rect 3644 4456 3652 4464
rect 2412 4436 2420 4444
rect 4076 4436 4084 4444
rect 4220 4436 4228 4444
rect 4412 4436 4420 4444
rect 5052 4436 5060 4444
rect 5468 4436 5476 4444
rect 5612 4436 5620 4444
rect 5740 4436 5748 4444
rect 6124 4436 6132 4444
rect 1577 4406 1585 4414
rect 1587 4406 1595 4414
rect 1597 4406 1605 4414
rect 1607 4406 1615 4414
rect 4665 4406 4673 4414
rect 4675 4406 4683 4414
rect 4685 4406 4693 4414
rect 4695 4406 4703 4414
rect 588 4376 596 4384
rect 892 4376 900 4384
rect 972 4376 980 4384
rect 1164 4376 1172 4384
rect 1404 4376 1412 4384
rect 1420 4376 1428 4384
rect 1580 4376 1588 4384
rect 1676 4376 1684 4384
rect 2284 4376 2292 4384
rect 2652 4376 2660 4384
rect 2812 4376 2820 4384
rect 2892 4376 2900 4384
rect 2956 4376 2964 4384
rect 3532 4376 3540 4384
rect 4332 4376 4340 4384
rect 4428 4376 4436 4384
rect 5788 4376 5796 4384
rect 6028 4376 6036 4384
rect 6156 4376 6164 4384
rect 12 4356 20 4364
rect 3772 4356 3780 4364
rect 5916 4356 5924 4364
rect 6204 4356 6212 4364
rect 1036 4336 1044 4344
rect 2204 4336 2212 4344
rect 2636 4336 2644 4344
rect 3356 4336 3364 4344
rect 4188 4336 4196 4344
rect 5628 4336 5636 4344
rect 940 4316 948 4324
rect 1004 4316 1012 4324
rect 1532 4316 1540 4324
rect 2236 4316 2244 4324
rect 140 4294 148 4302
rect 300 4296 308 4304
rect 476 4296 484 4304
rect 620 4296 628 4304
rect 700 4296 708 4304
rect 732 4296 740 4304
rect 828 4296 836 4304
rect 924 4296 932 4304
rect 1004 4296 1012 4304
rect 1036 4296 1044 4304
rect 1260 4296 1268 4304
rect 1372 4296 1380 4304
rect 1500 4296 1508 4304
rect 1548 4296 1556 4304
rect 1644 4296 1652 4304
rect 1772 4296 1780 4304
rect 1916 4296 1924 4304
rect 1932 4296 1940 4304
rect 1980 4296 1988 4304
rect 1996 4296 2004 4304
rect 2092 4296 2100 4304
rect 2124 4296 2132 4304
rect 2380 4316 2388 4324
rect 2428 4316 2436 4324
rect 3036 4316 3044 4324
rect 3608 4316 3616 4324
rect 2284 4296 2292 4304
rect 2540 4296 2548 4304
rect 2556 4296 2564 4304
rect 2684 4296 2692 4304
rect 2700 4296 2708 4304
rect 2732 4296 2740 4304
rect 2748 4296 2756 4304
rect 2780 4296 2788 4304
rect 2828 4296 2836 4304
rect 2844 4296 2852 4304
rect 2860 4296 2868 4304
rect 2924 4296 2932 4304
rect 2972 4296 2980 4304
rect 2988 4296 2996 4304
rect 3004 4296 3012 4304
rect 3228 4296 3236 4304
rect 3276 4296 3284 4304
rect 3372 4296 3380 4304
rect 3388 4296 3396 4304
rect 3404 4296 3412 4304
rect 3500 4296 3508 4304
rect 3548 4296 3556 4304
rect 3564 4296 3572 4304
rect 3596 4296 3604 4304
rect 3644 4316 3652 4324
rect 3756 4316 3764 4324
rect 3964 4316 3972 4324
rect 4204 4316 4212 4324
rect 4508 4316 4516 4324
rect 3884 4296 3892 4304
rect 4060 4294 4068 4302
rect 4284 4296 4292 4304
rect 4300 4296 4308 4304
rect 4348 4296 4356 4304
rect 4380 4296 4388 4304
rect 4396 4296 4404 4304
rect 4444 4296 4452 4304
rect 4652 4316 4660 4324
rect 4700 4316 4708 4324
rect 5164 4316 5172 4324
rect 4556 4296 4564 4304
rect 4604 4296 4612 4304
rect 4860 4296 4868 4304
rect 5384 4316 5392 4324
rect 5404 4316 5412 4324
rect 5692 4316 5700 4324
rect 5756 4316 5764 4324
rect 5820 4316 5828 4324
rect 5840 4316 5848 4324
rect 5884 4316 5892 4324
rect 6124 4316 6132 4324
rect 5068 4294 5076 4302
rect 5228 4296 5236 4304
rect 5372 4296 5380 4304
rect 5452 4296 5460 4304
rect 5516 4296 5524 4304
rect 5580 4296 5588 4304
rect 5612 4296 5620 4304
rect 5660 4296 5668 4304
rect 5756 4296 5764 4304
rect 5788 4296 5796 4304
rect 5852 4296 5860 4304
rect 5916 4296 5924 4304
rect 5948 4296 5956 4304
rect 6172 4296 6180 4304
rect 6220 4296 6228 4304
rect 268 4276 276 4284
rect 460 4276 468 4284
rect 508 4276 516 4284
rect 860 4276 868 4284
rect 1068 4276 1076 4284
rect 1084 4276 1092 4284
rect 1244 4276 1252 4284
rect 1452 4276 1460 4284
rect 876 4256 884 4264
rect 1068 4256 1076 4264
rect 1484 4276 1492 4284
rect 1820 4276 1828 4284
rect 1916 4276 1924 4284
rect 2204 4276 2212 4284
rect 2300 4276 2308 4284
rect 2396 4276 2404 4284
rect 2428 4276 2436 4284
rect 3580 4276 3588 4284
rect 3692 4276 3700 4284
rect 3900 4276 3908 4284
rect 3996 4276 4004 4284
rect 4076 4276 4084 4284
rect 4204 4276 4212 4284
rect 4252 4276 4260 4284
rect 4268 4276 4276 4284
rect 4460 4276 4468 4284
rect 4588 4276 4596 4284
rect 4652 4276 4660 4284
rect 4732 4276 4740 4284
rect 4908 4276 4916 4284
rect 5052 4276 5060 4284
rect 5180 4276 5188 4284
rect 5228 4276 5236 4284
rect 5244 4276 5252 4284
rect 5340 4276 5348 4284
rect 5356 4276 5364 4284
rect 5420 4276 5428 4284
rect 5468 4276 5476 4284
rect 5532 4276 5540 4284
rect 5564 4276 5572 4284
rect 5740 4276 5748 4284
rect 5804 4276 5812 4284
rect 5868 4276 5876 4284
rect 5932 4276 5940 4284
rect 5980 4276 5988 4284
rect 6060 4276 6068 4284
rect 6092 4276 6100 4284
rect 6172 4276 6180 4284
rect 6220 4276 6228 4284
rect 1532 4256 1540 4264
rect 1884 4256 1892 4264
rect 2316 4256 2324 4264
rect 2636 4256 2644 4264
rect 3020 4256 3028 4264
rect 3116 4256 3124 4264
rect 3356 4256 3364 4264
rect 3420 4256 3428 4264
rect 4252 4256 4260 4264
rect 4652 4256 4660 4264
rect 5436 4256 5444 4264
rect 5500 4256 5508 4264
rect 5980 4256 5988 4264
rect 6012 4256 6020 4264
rect 6044 4256 6052 4264
rect 6188 4256 6196 4264
rect 6268 4256 6276 4264
rect 572 4236 580 4244
rect 812 4236 820 4244
rect 1356 4236 1364 4244
rect 1692 4236 1700 4244
rect 2380 4236 2388 4244
rect 2412 4236 2420 4244
rect 3052 4236 3060 4244
rect 3740 4236 3748 4244
rect 3980 4236 3988 4244
rect 4524 4236 4532 4244
rect 4748 4236 4756 4244
rect 5276 4236 5284 4244
rect 5484 4236 5492 4244
rect 5548 4236 5556 4244
rect 3113 4206 3121 4214
rect 3123 4206 3131 4214
rect 3133 4206 3141 4214
rect 3143 4206 3151 4214
rect 188 4176 196 4184
rect 204 4176 212 4184
rect 860 4176 868 4184
rect 956 4176 964 4184
rect 1100 4176 1108 4184
rect 1340 4176 1348 4184
rect 1372 4176 1380 4184
rect 1404 4176 1412 4184
rect 1468 4176 1476 4184
rect 1708 4176 1716 4184
rect 1836 4176 1844 4184
rect 2044 4176 2052 4184
rect 2940 4176 2948 4184
rect 2988 4176 2996 4184
rect 3212 4176 3220 4184
rect 3292 4176 3300 4184
rect 3324 4176 3332 4184
rect 3548 4176 3556 4184
rect 3628 4176 3636 4184
rect 3772 4176 3780 4184
rect 3788 4176 3796 4184
rect 3996 4176 4004 4184
rect 4060 4176 4068 4184
rect 4396 4176 4404 4184
rect 4428 4176 4436 4184
rect 4620 4176 4628 4184
rect 4828 4176 4836 4184
rect 5724 4176 5732 4184
rect 5948 4176 5956 4184
rect 6076 4176 6084 4184
rect 284 4156 292 4164
rect 332 4156 340 4164
rect 508 4156 516 4164
rect 652 4156 660 4164
rect 732 4156 740 4164
rect 876 4156 884 4164
rect 892 4156 900 4164
rect 1324 4156 1332 4164
rect 1452 4156 1460 4164
rect 1596 4156 1604 4164
rect 1756 4156 1764 4164
rect 2028 4156 2036 4164
rect 2172 4156 2180 4164
rect 2428 4156 2436 4164
rect 2492 4156 2500 4164
rect 2828 4156 2836 4164
rect 3148 4156 3156 4164
rect 3308 4156 3316 4164
rect 3420 4156 3428 4164
rect 3564 4156 3572 4164
rect 348 4136 356 4144
rect 412 4136 420 4144
rect 428 4136 436 4144
rect 668 4136 676 4144
rect 908 4136 916 4144
rect 972 4136 980 4144
rect 1036 4136 1044 4144
rect 1324 4136 1332 4144
rect 1388 4136 1396 4144
rect 1436 4136 1444 4144
rect 1516 4136 1524 4144
rect 1692 4136 1700 4144
rect 1740 4136 1748 4144
rect 1772 4136 1780 4144
rect 1932 4136 1940 4144
rect 2492 4136 2500 4144
rect 2556 4136 2564 4144
rect 2860 4136 2868 4144
rect 3228 4136 3236 4144
rect 3340 4136 3348 4144
rect 76 4116 84 4124
rect 124 4116 132 4124
rect 236 4116 244 4124
rect 284 4116 292 4124
rect 364 4116 372 4124
rect 508 4118 516 4126
rect 748 4116 756 4124
rect 908 4116 916 4124
rect 972 4116 980 4124
rect 1052 4116 1060 4124
rect 204 4096 212 4104
rect 956 4096 964 4104
rect 988 4096 996 4104
rect 1020 4096 1028 4104
rect 1084 4096 1092 4104
rect 1148 4116 1156 4124
rect 1244 4116 1252 4124
rect 1308 4116 1316 4124
rect 1500 4116 1508 4124
rect 1580 4116 1588 4124
rect 1596 4116 1604 4124
rect 1644 4116 1652 4124
rect 1676 4116 1684 4124
rect 1788 4116 1796 4124
rect 1868 4116 1876 4124
rect 1884 4116 1892 4124
rect 1980 4116 1988 4124
rect 2156 4116 2164 4124
rect 2284 4116 2292 4124
rect 2412 4116 2420 4124
rect 1260 4096 1268 4104
rect 1292 4096 1300 4104
rect 1356 4096 1364 4104
rect 1468 4096 1476 4104
rect 1548 4096 1556 4104
rect 1644 4096 1652 4104
rect 1820 4096 1828 4104
rect 1948 4096 1956 4104
rect 1980 4096 1988 4104
rect 2604 4116 2612 4124
rect 2668 4116 2676 4124
rect 2716 4116 2724 4124
rect 2780 4116 2788 4124
rect 2828 4116 2836 4124
rect 2876 4116 2884 4124
rect 2908 4116 2916 4124
rect 2972 4116 2980 4124
rect 3052 4116 3060 4124
rect 3100 4116 3108 4124
rect 3244 4116 3252 4124
rect 3260 4116 3268 4124
rect 3356 4116 3364 4124
rect 3436 4116 3444 4124
rect 3564 4116 3572 4124
rect 3596 4116 3604 4124
rect 3612 4116 3620 4124
rect 3660 4116 3668 4124
rect 3708 4116 3716 4124
rect 4124 4156 4132 4164
rect 4172 4156 4180 4164
rect 4412 4156 4420 4164
rect 4684 4156 4692 4164
rect 4812 4156 4820 4164
rect 4956 4156 4964 4164
rect 5084 4156 5092 4164
rect 5436 4156 5444 4164
rect 5468 4156 5476 4164
rect 4444 4136 4452 4144
rect 4540 4136 4548 4144
rect 4780 4136 4788 4144
rect 5084 4136 5092 4144
rect 5116 4136 5124 4144
rect 5228 4136 5236 4144
rect 5260 4136 5268 4144
rect 5340 4136 5348 4144
rect 5404 4136 5412 4144
rect 5484 4136 5492 4144
rect 5516 4136 5524 4144
rect 5564 4136 5572 4144
rect 5660 4136 5668 4144
rect 5676 4136 5684 4144
rect 5788 4136 5796 4144
rect 5916 4136 5924 4144
rect 5932 4136 5940 4144
rect 6044 4136 6052 4144
rect 6060 4136 6068 4144
rect 6124 4136 6132 4144
rect 6188 4136 6196 4144
rect 3836 4116 3844 4124
rect 3916 4116 3924 4124
rect 3964 4116 3972 4124
rect 4012 4116 4020 4124
rect 4028 4116 4036 4124
rect 4076 4116 4084 4124
rect 4092 4116 4100 4124
rect 4156 4116 4164 4124
rect 4204 4116 4212 4124
rect 4236 4116 4244 4124
rect 4300 4116 4308 4124
rect 4364 4116 4372 4124
rect 4524 4116 4532 4124
rect 4700 4116 4708 4124
rect 4716 4116 4724 4124
rect 4764 4116 4772 4124
rect 4940 4116 4948 4124
rect 5020 4116 5028 4124
rect 5052 4116 5060 4124
rect 5100 4116 5108 4124
rect 5180 4116 5188 4124
rect 5244 4116 5252 4124
rect 2556 4096 2564 4104
rect 2620 4096 2628 4104
rect 2684 4096 2692 4104
rect 2700 4096 2708 4104
rect 2764 4096 2772 4104
rect 2892 4096 2900 4104
rect 2956 4096 2964 4104
rect 3020 4096 3028 4104
rect 3084 4096 3092 4104
rect 3692 4096 3700 4104
rect 3756 4096 3764 4104
rect 3820 4096 3828 4104
rect 3932 4096 3940 4104
rect 3948 4096 3956 4104
rect 4156 4096 4164 4104
rect 4252 4096 4260 4104
rect 4316 4096 4324 4104
rect 4332 4096 4340 4104
rect 4380 4096 4388 4104
rect 4748 4096 4756 4104
rect 5020 4096 5028 4104
rect 5148 4096 5156 4104
rect 5212 4096 5220 4104
rect 5324 4116 5332 4124
rect 5372 4116 5380 4124
rect 5388 4116 5396 4124
rect 5500 4116 5508 4124
rect 5292 4096 5300 4104
rect 5324 4096 5332 4104
rect 5356 4096 5364 4104
rect 5548 4116 5556 4124
rect 5676 4116 5684 4124
rect 5772 4116 5780 4124
rect 5740 4096 5748 4104
rect 5852 4096 5860 4104
rect 5916 4116 5924 4124
rect 5980 4116 5988 4124
rect 6028 4116 6036 4124
rect 6060 4116 6068 4124
rect 6124 4116 6132 4124
rect 6140 4116 6148 4124
rect 6188 4116 6196 4124
rect 6220 4116 6228 4124
rect 5996 4096 6004 4104
rect 6140 4096 6148 4104
rect 6172 4096 6180 4104
rect 6220 4096 6228 4104
rect 316 4076 324 4084
rect 636 4076 644 4084
rect 2492 4076 2500 4084
rect 2588 4076 2596 4084
rect 2620 4076 2628 4084
rect 2652 4076 2660 4084
rect 2668 4076 2676 4084
rect 364 4056 372 4064
rect 1212 4056 1220 4064
rect 2732 4076 2740 4084
rect 2796 4076 2804 4084
rect 2924 4076 2932 4084
rect 2956 4076 2964 4084
rect 3052 4076 3060 4084
rect 3116 4076 3124 4084
rect 3724 4076 3732 4084
rect 3788 4076 3796 4084
rect 3852 4076 3860 4084
rect 3900 4076 3908 4084
rect 3980 4076 3988 4084
rect 4172 4076 4180 4084
rect 4220 4076 4228 4084
rect 4268 4076 4276 4084
rect 4284 4076 4292 4084
rect 4348 4076 4356 4084
rect 6236 4076 6244 4084
rect 3036 4056 3044 4064
rect 3100 4056 3108 4064
rect 3836 4056 3844 4064
rect 5420 4056 5428 4064
rect 892 4036 900 4044
rect 1164 4036 1172 4044
rect 1340 4036 1348 4044
rect 1788 4036 1796 4044
rect 2012 4036 2020 4044
rect 2300 4036 2308 4044
rect 2604 4036 2612 4044
rect 2780 4036 2788 4044
rect 2908 4036 2916 4044
rect 3148 4036 3156 4044
rect 3180 4036 3188 4044
rect 3708 4036 3716 4044
rect 3884 4036 3892 4044
rect 5180 4036 5188 4044
rect 5900 4036 5908 4044
rect 6220 4036 6228 4044
rect 1577 4006 1585 4014
rect 1587 4006 1595 4014
rect 1597 4006 1605 4014
rect 1607 4006 1615 4014
rect 4665 4006 4673 4014
rect 4675 4006 4683 4014
rect 4685 4006 4693 4014
rect 4695 4006 4703 4014
rect 172 3976 180 3984
rect 492 3976 500 3984
rect 556 3976 564 3984
rect 1356 3976 1364 3984
rect 1804 3976 1812 3984
rect 1900 3976 1908 3984
rect 2156 3976 2164 3984
rect 2236 3976 2244 3984
rect 2252 3976 2260 3984
rect 2460 3976 2468 3984
rect 2508 3976 2516 3984
rect 2524 3976 2532 3984
rect 2860 3976 2868 3984
rect 2876 3976 2884 3984
rect 3292 3976 3300 3984
rect 3596 3976 3604 3984
rect 3644 3976 3652 3984
rect 3692 3976 3700 3984
rect 3900 3976 3908 3984
rect 4076 3976 4084 3984
rect 4636 3976 4644 3984
rect 5852 3976 5860 3984
rect 5948 3976 5956 3984
rect 76 3956 84 3964
rect 2796 3956 2804 3964
rect 3484 3956 3492 3964
rect 6076 3956 6084 3964
rect 252 3936 260 3944
rect 812 3936 820 3944
rect 1276 3936 1284 3944
rect 1772 3936 1780 3944
rect 2332 3936 2340 3944
rect 2364 3936 2372 3944
rect 2780 3936 2788 3944
rect 3420 3936 3428 3944
rect 3500 3936 3508 3944
rect 3564 3936 3572 3944
rect 3708 3936 3716 3944
rect 3788 3936 3796 3944
rect 3980 3936 3988 3944
rect 92 3916 100 3924
rect 380 3916 388 3924
rect 412 3916 420 3924
rect 444 3916 452 3924
rect 460 3916 468 3924
rect 860 3916 868 3924
rect 76 3896 84 3904
rect 124 3896 132 3904
rect 172 3896 180 3904
rect 268 3896 276 3904
rect 348 3896 356 3904
rect 412 3896 420 3904
rect 524 3896 532 3904
rect 684 3896 692 3904
rect 860 3896 868 3904
rect 908 3916 916 3924
rect 1100 3916 1108 3924
rect 1132 3916 1140 3924
rect 1260 3916 1268 3924
rect 1388 3916 1396 3924
rect 1452 3916 1460 3924
rect 1532 3916 1540 3924
rect 1692 3916 1700 3924
rect 1884 3916 1892 3924
rect 1964 3916 1972 3924
rect 2028 3916 2036 3924
rect 2140 3916 2148 3924
rect 2396 3916 2404 3924
rect 2716 3916 2724 3924
rect 2748 3916 2756 3924
rect 2812 3916 2820 3924
rect 1020 3896 1028 3904
rect 1132 3896 1140 3904
rect 1148 3896 1156 3904
rect 1484 3896 1492 3904
rect 1548 3896 1556 3904
rect 1724 3896 1732 3904
rect 1820 3896 1828 3904
rect 108 3876 116 3884
rect 140 3876 148 3884
rect 156 3876 164 3884
rect 220 3876 228 3884
rect 236 3876 244 3884
rect 284 3876 292 3884
rect 332 3876 340 3884
rect 364 3876 372 3884
rect 508 3876 516 3884
rect 572 3876 580 3884
rect 604 3876 612 3884
rect 636 3876 644 3884
rect 844 3876 852 3884
rect 940 3876 948 3884
rect 1036 3876 1044 3884
rect 1084 3876 1092 3884
rect 1148 3876 1156 3884
rect 1212 3876 1220 3884
rect 1404 3876 1412 3884
rect 1516 3876 1524 3884
rect 1580 3876 1588 3884
rect 1644 3876 1652 3884
rect 1820 3876 1828 3884
rect 1996 3896 2004 3904
rect 2188 3896 2196 3904
rect 2204 3896 2212 3904
rect 2380 3896 2388 3904
rect 2428 3896 2436 3904
rect 2476 3896 2484 3904
rect 2604 3896 2612 3904
rect 2780 3896 2788 3904
rect 2860 3896 2868 3904
rect 2940 3896 2948 3904
rect 3036 3896 3044 3904
rect 3164 3916 3172 3924
rect 3468 3916 3476 3924
rect 3532 3916 3540 3924
rect 3740 3916 3748 3924
rect 3756 3916 3764 3924
rect 3820 3916 3828 3924
rect 3948 3916 3956 3924
rect 4012 3916 4020 3924
rect 3180 3896 3188 3904
rect 3260 3896 3268 3904
rect 3324 3896 3332 3904
rect 3372 3896 3380 3904
rect 3452 3896 3460 3904
rect 3484 3896 3492 3904
rect 3548 3896 3556 3904
rect 3628 3896 3636 3904
rect 3676 3896 3684 3904
rect 3724 3896 3732 3904
rect 3772 3896 3780 3904
rect 3932 3896 3940 3904
rect 3980 3896 3988 3904
rect 1964 3876 1972 3884
rect 2044 3876 2052 3884
rect 2092 3876 2100 3884
rect 2108 3876 2116 3884
rect 2284 3876 2292 3884
rect 2556 3876 2564 3884
rect 2588 3876 2596 3884
rect 2652 3876 2660 3884
rect 2668 3880 2676 3888
rect 2716 3876 2724 3884
rect 2924 3876 2932 3884
rect 2988 3876 2996 3884
rect 3148 3876 3156 3884
rect 3164 3876 3172 3884
rect 3276 3876 3284 3884
rect 3388 3876 3396 3884
rect 4076 3936 4084 3944
rect 4092 3936 4100 3944
rect 4204 3936 4212 3944
rect 4236 3936 4244 3944
rect 5020 3936 5028 3944
rect 5772 3936 5780 3944
rect 5996 3936 6004 3944
rect 4060 3916 4068 3924
rect 4076 3916 4084 3924
rect 4124 3916 4132 3924
rect 4220 3916 4228 3924
rect 4268 3916 4276 3924
rect 4124 3896 4132 3904
rect 4172 3896 4180 3904
rect 4252 3896 4260 3904
rect 4284 3896 4292 3904
rect 4348 3916 4356 3924
rect 5052 3916 5060 3924
rect 5068 3916 5076 3924
rect 5132 3916 5140 3924
rect 5404 3916 5412 3924
rect 5436 3916 5444 3924
rect 5628 3916 5636 3924
rect 5660 3916 5668 3924
rect 5676 3916 5684 3924
rect 5740 3916 5748 3924
rect 5980 3916 5988 3924
rect 6252 3916 6260 3924
rect 4508 3896 4516 3904
rect 4764 3894 4772 3902
rect 4956 3894 4964 3902
rect 5164 3896 5172 3904
rect 5196 3896 5204 3904
rect 5340 3896 5348 3904
rect 5404 3896 5412 3904
rect 5468 3896 5476 3904
rect 5484 3896 5492 3904
rect 5708 3896 5716 3904
rect 5772 3896 5780 3904
rect 5788 3896 5796 3904
rect 5820 3896 5828 3904
rect 5884 3896 5892 3904
rect 5916 3896 5924 3904
rect 6028 3896 6036 3904
rect 6060 3896 6068 3904
rect 6124 3896 6132 3904
rect 6156 3896 6164 3904
rect 6188 3896 6196 3904
rect 6236 3896 6244 3904
rect 4156 3876 4164 3884
rect 4284 3876 4292 3884
rect 4348 3876 4356 3884
rect 4508 3876 4516 3884
rect 4556 3876 4564 3884
rect 4796 3876 4804 3884
rect 4940 3876 4948 3884
rect 5052 3876 5060 3884
rect 5116 3876 5124 3884
rect 5180 3876 5188 3884
rect 5196 3876 5204 3884
rect 12 3856 20 3864
rect 44 3856 52 3864
rect 316 3856 324 3864
rect 668 3856 676 3864
rect 812 3856 820 3864
rect 956 3856 964 3864
rect 1068 3856 1076 3864
rect 1196 3856 1204 3864
rect 2092 3856 2100 3864
rect 2252 3856 2260 3864
rect 2316 3856 2324 3864
rect 2524 3856 2532 3864
rect 2828 3856 2836 3864
rect 2908 3856 2916 3864
rect 3052 3856 3060 3864
rect 3884 3856 3892 3864
rect 4012 3856 4020 3864
rect 4700 3856 4708 3864
rect 5292 3876 5300 3884
rect 5324 3876 5332 3884
rect 5372 3876 5380 3884
rect 5500 3876 5508 3884
rect 5532 3876 5540 3884
rect 5596 3876 5604 3884
rect 5660 3876 5668 3884
rect 5724 3876 5732 3884
rect 5788 3876 5796 3884
rect 5836 3876 5844 3884
rect 5868 3876 5876 3884
rect 5932 3876 5940 3884
rect 5996 3876 6004 3884
rect 6044 3876 6052 3884
rect 6076 3876 6084 3884
rect 6140 3876 6148 3884
rect 6172 3876 6180 3884
rect 6204 3876 6212 3884
rect 5244 3856 5252 3864
rect 5372 3856 5380 3864
rect 5452 3856 5460 3864
rect 5612 3856 5620 3864
rect 5628 3856 5636 3864
rect 5836 3856 5844 3864
rect 5916 3856 5924 3864
rect 6140 3856 6148 3864
rect 300 3836 308 3844
rect 972 3836 980 3844
rect 1052 3836 1060 3844
rect 1180 3836 1188 3844
rect 2364 3836 2372 3844
rect 2636 3836 2644 3844
rect 2732 3836 2740 3844
rect 2972 3836 2980 3844
rect 3068 3836 3076 3844
rect 3212 3836 3220 3844
rect 3340 3836 3348 3844
rect 3580 3836 3588 3844
rect 3772 3836 3780 3844
rect 3836 3836 3844 3844
rect 4396 3836 4404 3844
rect 5308 3836 5316 3844
rect 5356 3836 5364 3844
rect 5516 3836 5524 3844
rect 5852 3836 5860 3844
rect 5900 3836 5908 3844
rect 3113 3806 3121 3814
rect 3123 3806 3131 3814
rect 3133 3806 3141 3814
rect 3143 3806 3151 3814
rect 156 3776 164 3784
rect 332 3776 340 3784
rect 460 3776 468 3784
rect 636 3776 644 3784
rect 828 3776 836 3784
rect 844 3776 852 3784
rect 908 3776 916 3784
rect 1164 3776 1172 3784
rect 1484 3776 1492 3784
rect 1564 3776 1572 3784
rect 1900 3776 1908 3784
rect 2348 3776 2356 3784
rect 2412 3776 2420 3784
rect 2428 3776 2436 3784
rect 2796 3776 2804 3784
rect 3084 3776 3092 3784
rect 3260 3776 3268 3784
rect 3388 3776 3396 3784
rect 3612 3776 3620 3784
rect 3788 3776 3796 3784
rect 3852 3776 3860 3784
rect 4172 3776 4180 3784
rect 4348 3776 4356 3784
rect 60 3756 68 3764
rect 236 3756 244 3764
rect 924 3756 932 3764
rect 1036 3756 1044 3764
rect 1116 3756 1124 3764
rect 1260 3756 1268 3764
rect 44 3736 52 3744
rect 76 3736 84 3744
rect 140 3736 148 3744
rect 204 3736 212 3744
rect 316 3736 324 3744
rect 364 3736 372 3744
rect 412 3736 420 3744
rect 444 3736 452 3744
rect 460 3736 468 3744
rect 492 3736 500 3744
rect 540 3736 548 3744
rect 588 3736 596 3744
rect 668 3736 676 3744
rect 860 3736 868 3744
rect 876 3736 884 3744
rect 988 3736 996 3744
rect 1052 3736 1060 3744
rect 1084 3736 1092 3744
rect 1116 3736 1124 3744
rect 1212 3736 1220 3744
rect 1276 3736 1284 3744
rect 1308 3736 1316 3744
rect 1372 3736 1380 3744
rect 1420 3736 1428 3744
rect 2028 3756 2036 3764
rect 3020 3756 3028 3764
rect 3372 3756 3380 3764
rect 3676 3756 3684 3764
rect 3740 3756 3748 3764
rect 3964 3756 3972 3764
rect 4332 3756 4340 3764
rect 4940 3776 4948 3784
rect 4988 3776 4996 3784
rect 5196 3776 5204 3784
rect 5260 3776 5268 3784
rect 5676 3776 5684 3784
rect 5740 3776 5748 3784
rect 5884 3776 5892 3784
rect 5996 3776 6004 3784
rect 6044 3776 6052 3784
rect 6092 3776 6100 3784
rect 6252 3776 6260 3784
rect 5164 3756 5172 3764
rect 5436 3756 5444 3764
rect 5484 3756 5492 3764
rect 5660 3756 5668 3764
rect 5724 3756 5732 3764
rect 6188 3756 6196 3764
rect 1468 3736 1476 3744
rect 1484 3736 1492 3744
rect 1564 3736 1572 3744
rect 1804 3736 1812 3744
rect 1820 3736 1828 3744
rect 1884 3736 1892 3744
rect 1996 3736 2004 3744
rect 92 3716 100 3724
rect 140 3716 148 3724
rect 172 3716 180 3724
rect 268 3716 276 3724
rect 300 3716 308 3724
rect 412 3716 420 3724
rect 444 3716 452 3724
rect 508 3716 516 3724
rect 540 3716 548 3724
rect 588 3716 596 3724
rect 700 3718 708 3726
rect 876 3716 884 3724
rect 988 3716 996 3724
rect 1004 3716 1012 3724
rect 1068 3716 1076 3724
rect 1148 3716 1156 3724
rect 1212 3716 1220 3724
rect 1228 3716 1236 3724
rect 1324 3716 1332 3724
rect 1388 3716 1396 3724
rect 1404 3716 1412 3724
rect 1468 3716 1476 3724
rect 1548 3716 1556 3724
rect 1660 3716 1668 3724
rect 1724 3716 1732 3724
rect 1804 3716 1812 3724
rect 1836 3716 1844 3724
rect 1884 3716 1892 3724
rect 2028 3716 2036 3724
rect 2060 3716 2068 3724
rect 2124 3736 2132 3744
rect 2156 3736 2164 3744
rect 2364 3736 2372 3744
rect 2780 3736 2788 3744
rect 2812 3736 2820 3744
rect 2828 3736 2836 3744
rect 3308 3736 3316 3744
rect 3404 3736 3412 3744
rect 3628 3736 3636 3744
rect 3724 3736 3732 3744
rect 3868 3736 3876 3744
rect 4204 3736 4212 3744
rect 4284 3736 4292 3744
rect 4300 3736 4308 3744
rect 4476 3736 4484 3744
rect 4508 3736 4516 3744
rect 4636 3736 4644 3744
rect 4876 3736 4884 3744
rect 4972 3736 4980 3744
rect 5084 3736 5092 3744
rect 5100 3736 5108 3744
rect 5180 3736 5188 3744
rect 5244 3736 5252 3744
rect 5372 3736 5380 3744
rect 5388 3736 5396 3744
rect 5452 3736 5460 3744
rect 5468 3736 5476 3744
rect 5532 3736 5540 3744
rect 5628 3736 5636 3744
rect 5724 3736 5732 3744
rect 5756 3736 5764 3744
rect 5772 3736 5780 3744
rect 5820 3736 5828 3744
rect 5836 3736 5844 3744
rect 5900 3736 5908 3744
rect 5916 3736 5924 3744
rect 5964 3736 5972 3744
rect 6012 3736 6020 3744
rect 6060 3736 6068 3744
rect 6108 3736 6116 3744
rect 6188 3736 6196 3744
rect 6252 3736 6260 3744
rect 6284 3736 6292 3744
rect 140 3696 148 3704
rect 172 3696 180 3704
rect 332 3696 340 3704
rect 412 3696 420 3704
rect 524 3696 532 3704
rect 636 3696 644 3704
rect 940 3696 948 3704
rect 1100 3696 1108 3704
rect 1164 3696 1172 3704
rect 1324 3696 1332 3704
rect 1724 3696 1732 3704
rect 2012 3696 2020 3704
rect 2252 3716 2260 3724
rect 2460 3716 2468 3724
rect 2556 3716 2564 3724
rect 2684 3716 2692 3724
rect 2700 3716 2708 3724
rect 2764 3716 2772 3724
rect 2412 3696 2420 3704
rect 2428 3696 2436 3704
rect 2860 3716 2868 3724
rect 2908 3716 2916 3724
rect 2924 3716 2932 3724
rect 2972 3716 2980 3724
rect 3196 3716 3204 3724
rect 3228 3716 3236 3724
rect 3340 3716 3348 3724
rect 3356 3716 3364 3724
rect 3420 3716 3428 3724
rect 3516 3716 3524 3724
rect 2812 3696 2820 3704
rect 2892 3696 2900 3704
rect 3004 3696 3012 3704
rect 3084 3696 3092 3704
rect 3164 3696 3172 3704
rect 3228 3696 3236 3704
rect 3308 3696 3316 3704
rect 3660 3696 3668 3704
rect 3708 3716 3716 3724
rect 3820 3716 3828 3724
rect 3916 3716 3924 3724
rect 3932 3716 3940 3724
rect 3996 3716 4004 3724
rect 4076 3716 4084 3724
rect 4140 3716 4148 3724
rect 4220 3716 4228 3724
rect 4236 3716 4244 3724
rect 4300 3716 4308 3724
rect 4460 3716 4468 3724
rect 4540 3716 4548 3724
rect 4556 3716 4564 3724
rect 4604 3716 4612 3724
rect 4828 3716 4836 3724
rect 4908 3716 4916 3724
rect 5036 3716 5044 3724
rect 5148 3716 5156 3724
rect 5228 3716 5236 3724
rect 5292 3716 5300 3724
rect 5356 3716 5364 3724
rect 5388 3716 5396 3724
rect 5532 3716 5540 3724
rect 5580 3716 5588 3724
rect 5756 3716 5764 3724
rect 5788 3716 5796 3724
rect 5820 3716 5828 3724
rect 5852 3716 5860 3724
rect 5884 3716 5892 3724
rect 5932 3716 5940 3724
rect 6124 3716 6132 3724
rect 6140 3716 6148 3724
rect 3804 3696 3812 3704
rect 3980 3696 3988 3704
rect 4092 3696 4100 3704
rect 4156 3696 4164 3704
rect 4172 3696 4180 3704
rect 4588 3696 4596 3704
rect 5004 3696 5012 3704
rect 5116 3696 5124 3704
rect 5196 3696 5204 3704
rect 5324 3696 5332 3704
rect 5436 3696 5444 3704
rect 5516 3696 5524 3704
rect 5580 3696 5588 3704
rect 5676 3696 5684 3704
rect 5948 3696 5956 3704
rect 5996 3696 6004 3704
rect 6044 3696 6052 3704
rect 6092 3696 6100 3704
rect 6156 3696 6164 3704
rect 6172 3696 6180 3704
rect 6236 3696 6244 3704
rect 6252 3696 6260 3704
rect 396 3676 404 3684
rect 556 3676 564 3684
rect 1004 3676 1012 3684
rect 1228 3676 1236 3684
rect 1452 3676 1460 3684
rect 2668 3676 2676 3684
rect 3980 3676 3988 3684
rect 300 3656 308 3664
rect 4012 3676 4020 3684
rect 4044 3676 4052 3684
rect 4060 3676 4068 3684
rect 4124 3676 4132 3684
rect 5548 3676 5556 3684
rect 5724 3676 5732 3684
rect 12 3636 20 3644
rect 972 3636 980 3644
rect 2092 3636 2100 3644
rect 4140 3636 4148 3644
rect 4668 3636 4676 3644
rect 4700 3636 4708 3644
rect 5452 3636 5460 3644
rect 5500 3636 5508 3644
rect 5644 3636 5652 3644
rect 1577 3606 1585 3614
rect 1587 3606 1595 3614
rect 1597 3606 1605 3614
rect 1607 3606 1615 3614
rect 4665 3606 4673 3614
rect 4675 3606 4683 3614
rect 4685 3606 4693 3614
rect 4695 3606 4703 3614
rect 172 3576 180 3584
rect 492 3576 500 3584
rect 572 3576 580 3584
rect 620 3576 628 3584
rect 748 3576 756 3584
rect 876 3576 884 3584
rect 1484 3576 1492 3584
rect 2108 3576 2116 3584
rect 2156 3576 2164 3584
rect 2188 3576 2196 3584
rect 2572 3576 2580 3584
rect 2700 3576 2708 3584
rect 2732 3576 2740 3584
rect 2908 3576 2916 3584
rect 3004 3576 3012 3584
rect 3084 3576 3092 3584
rect 3164 3576 3172 3584
rect 3324 3576 3332 3584
rect 3484 3576 3492 3584
rect 3788 3576 3796 3584
rect 3836 3576 3844 3584
rect 4716 3576 4724 3584
rect 5228 3576 5236 3584
rect 5356 3576 5364 3584
rect 5580 3576 5588 3584
rect 5756 3576 5764 3584
rect 5884 3576 5892 3584
rect 5980 3576 5988 3584
rect 6172 3576 6180 3584
rect 1180 3556 1188 3564
rect 1692 3556 1700 3564
rect 1884 3556 1892 3564
rect 2428 3556 2436 3564
rect 3564 3556 3572 3564
rect 6140 3556 6148 3564
rect 28 3536 36 3544
rect 556 3536 564 3544
rect 764 3536 772 3544
rect 908 3536 916 3544
rect 1116 3536 1124 3544
rect 1196 3536 1204 3544
rect 1468 3536 1476 3544
rect 2844 3536 2852 3544
rect 3228 3536 3236 3544
rect 3292 3536 3300 3544
rect 3692 3536 3700 3544
rect 3740 3536 3748 3544
rect 3980 3536 3988 3544
rect 4060 3536 4068 3544
rect 4140 3536 4148 3544
rect 4332 3536 4340 3544
rect 4732 3536 4740 3544
rect 4892 3536 4900 3544
rect 5372 3536 5380 3544
rect 5500 3536 5508 3544
rect 5900 3536 5908 3544
rect 60 3516 68 3524
rect 76 3516 84 3524
rect 524 3516 532 3524
rect 572 3516 580 3524
rect 796 3516 804 3524
rect 924 3516 932 3524
rect 988 3516 996 3524
rect 1164 3516 1172 3524
rect 1244 3516 1252 3524
rect 1276 3516 1284 3524
rect 1404 3516 1412 3524
rect 1468 3516 1476 3524
rect 1596 3516 1604 3524
rect 44 3496 52 3504
rect 76 3496 84 3504
rect 124 3496 132 3504
rect 172 3496 180 3504
rect 316 3496 324 3504
rect 428 3496 436 3504
rect 492 3496 500 3504
rect 572 3496 580 3504
rect 604 3496 612 3504
rect 668 3496 676 3504
rect 684 3496 692 3504
rect 780 3496 788 3504
rect 812 3496 820 3504
rect 892 3496 900 3504
rect 972 3496 980 3504
rect 1020 3496 1028 3504
rect 1036 3496 1044 3504
rect 1116 3496 1124 3504
rect 1180 3496 1188 3504
rect 1228 3496 1236 3504
rect 1292 3496 1300 3504
rect 1372 3496 1380 3504
rect 1420 3496 1428 3504
rect 1452 3496 1460 3504
rect 1484 3496 1492 3504
rect 1916 3516 1924 3524
rect 1948 3516 1956 3524
rect 2124 3516 2132 3524
rect 2460 3516 2468 3524
rect 3724 3516 3732 3524
rect 3964 3516 3972 3524
rect 4012 3516 4020 3524
rect 4092 3516 4100 3524
rect 4108 3516 4116 3524
rect 4172 3516 4180 3524
rect 4316 3516 4324 3524
rect 4556 3516 4564 3524
rect 1964 3496 1972 3504
rect 2060 3496 2068 3504
rect 2156 3496 2164 3504
rect 2332 3496 2340 3504
rect 2428 3496 2436 3504
rect 2524 3496 2532 3504
rect 2620 3496 2628 3504
rect 3100 3496 3108 3504
rect 3340 3496 3348 3504
rect 3388 3496 3396 3504
rect 3468 3496 3476 3504
rect 3756 3496 3764 3504
rect 3804 3496 3812 3504
rect 3852 3496 3860 3504
rect 3916 3496 3924 3504
rect 3932 3496 3940 3504
rect 3964 3496 3972 3504
rect 4076 3496 4084 3504
rect 4124 3496 4132 3504
rect 4220 3496 4228 3504
rect 4236 3496 4244 3504
rect 4300 3496 4308 3504
rect 4460 3496 4468 3504
rect 4556 3496 4564 3504
rect 4588 3496 4596 3504
rect 4636 3496 4644 3504
rect 4796 3496 4804 3504
rect 4844 3516 4852 3524
rect 5116 3516 5124 3524
rect 5180 3516 5188 3524
rect 5196 3516 5204 3524
rect 4972 3496 4980 3504
rect 5116 3496 5124 3504
rect 5228 3496 5236 3504
rect 5260 3496 5268 3504
rect 5324 3496 5332 3504
rect 5420 3496 5428 3504
rect 5484 3496 5492 3504
rect 5532 3496 5540 3504
rect 5564 3496 5572 3504
rect 5628 3516 5636 3524
rect 5660 3496 5668 3504
rect 5692 3496 5700 3504
rect 5804 3516 5812 3524
rect 5868 3516 5876 3524
rect 6204 3516 6212 3524
rect 5836 3496 5844 3504
rect 5884 3496 5892 3504
rect 6076 3496 6084 3504
rect 6188 3496 6196 3504
rect 44 3476 52 3484
rect 140 3476 148 3484
rect 188 3476 196 3484
rect 204 3480 212 3488
rect 332 3476 340 3484
rect 396 3476 404 3484
rect 412 3476 420 3484
rect 620 3476 628 3484
rect 652 3476 660 3484
rect 700 3476 708 3484
rect 828 3476 836 3484
rect 844 3476 852 3484
rect 972 3476 980 3484
rect 1036 3476 1044 3484
rect 1068 3476 1076 3484
rect 1228 3476 1236 3484
rect 1308 3476 1316 3484
rect 1436 3476 1444 3484
rect 1564 3476 1572 3484
rect 1596 3476 1604 3484
rect 1644 3476 1652 3484
rect 1660 3476 1668 3484
rect 1724 3476 1732 3484
rect 1756 3476 1764 3484
rect 1788 3476 1796 3484
rect 1836 3476 1844 3484
rect 1900 3476 1908 3484
rect 2028 3476 2036 3484
rect 2076 3476 2084 3484
rect 2172 3476 2180 3484
rect 2236 3476 2244 3484
rect 2540 3476 2548 3484
rect 2604 3476 2612 3484
rect 2796 3476 2804 3484
rect 2860 3476 2868 3484
rect 2876 3476 2884 3484
rect 2940 3476 2948 3484
rect 2956 3476 2964 3484
rect 3020 3476 3028 3484
rect 3036 3476 3044 3484
rect 3100 3476 3108 3484
rect 3164 3476 3172 3484
rect 3260 3476 3268 3484
rect 3420 3476 3428 3484
rect 3452 3476 3460 3484
rect 3516 3480 3524 3488
rect 3532 3476 3540 3484
rect 3548 3476 3556 3484
rect 3596 3476 3604 3484
rect 4204 3476 4212 3484
rect 4476 3476 4484 3484
rect 4780 3476 4788 3484
rect 4844 3476 4852 3484
rect 140 3456 148 3464
rect 348 3456 356 3464
rect 732 3456 740 3464
rect 860 3456 868 3464
rect 1100 3456 1108 3464
rect 1116 3456 1124 3464
rect 1148 3456 1156 3464
rect 1340 3456 1348 3464
rect 5084 3476 5092 3484
rect 5132 3476 5140 3484
rect 5180 3476 5188 3484
rect 5244 3476 5252 3484
rect 5276 3476 5284 3484
rect 5324 3476 5332 3484
rect 5420 3476 5428 3484
rect 5468 3476 5476 3484
rect 5548 3476 5556 3484
rect 5564 3476 5572 3484
rect 5596 3476 5604 3484
rect 5676 3476 5684 3484
rect 5740 3476 5748 3484
rect 5852 3476 5860 3484
rect 5964 3476 5972 3484
rect 6076 3476 6084 3484
rect 6236 3476 6244 3484
rect 1836 3456 1844 3464
rect 2028 3456 2036 3464
rect 2108 3456 2116 3464
rect 2204 3456 2212 3464
rect 2732 3456 2740 3464
rect 3148 3456 3156 3464
rect 3228 3456 3236 3464
rect 3420 3456 3428 3464
rect 4028 3456 4036 3464
rect 4332 3456 4340 3464
rect 4556 3456 4564 3464
rect 4732 3456 4740 3464
rect 4764 3456 4772 3464
rect 5020 3456 5028 3464
rect 5340 3456 5348 3464
rect 5404 3456 5412 3464
rect 5724 3456 5732 3464
rect 5932 3456 5940 3464
rect 6044 3456 6052 3464
rect 6076 3456 6084 3464
rect 6124 3456 6132 3464
rect 6156 3456 6164 3464
rect 6188 3456 6196 3464
rect 268 3436 276 3444
rect 332 3436 340 3444
rect 460 3436 468 3444
rect 716 3436 724 3444
rect 988 3436 996 3444
rect 1548 3436 1556 3444
rect 2668 3436 2676 3444
rect 3356 3436 3364 3444
rect 3644 3436 3652 3444
rect 3708 3436 3716 3444
rect 3884 3436 3892 3444
rect 3980 3436 3988 3444
rect 4044 3436 4052 3444
rect 4140 3436 4148 3444
rect 4172 3436 4180 3444
rect 4268 3436 4276 3444
rect 4620 3436 4628 3444
rect 5116 3436 5124 3444
rect 5292 3436 5300 3444
rect 5452 3436 5460 3444
rect 6060 3436 6068 3444
rect 3113 3406 3121 3414
rect 3123 3406 3131 3414
rect 3133 3406 3141 3414
rect 3143 3406 3151 3414
rect 188 3376 196 3384
rect 428 3376 436 3384
rect 940 3376 948 3384
rect 1228 3376 1236 3384
rect 1260 3376 1268 3384
rect 1484 3376 1492 3384
rect 1516 3376 1524 3384
rect 1900 3376 1908 3384
rect 2172 3376 2180 3384
rect 2332 3376 2340 3384
rect 2380 3376 2388 3384
rect 2572 3376 2580 3384
rect 3132 3376 3140 3384
rect 3164 3376 3172 3384
rect 3228 3376 3236 3384
rect 3596 3376 3604 3384
rect 3820 3376 3828 3384
rect 4044 3376 4052 3384
rect 4204 3376 4212 3384
rect 4348 3376 4356 3384
rect 4540 3376 4548 3384
rect 4892 3376 4900 3384
rect 5196 3376 5204 3384
rect 5276 3376 5284 3384
rect 556 3356 564 3364
rect 668 3356 676 3364
rect 1244 3356 1252 3364
rect 1420 3356 1428 3364
rect 2156 3356 2164 3364
rect 2396 3356 2404 3364
rect 76 3336 84 3344
rect 204 3336 212 3344
rect 508 3336 516 3344
rect 540 3336 548 3344
rect 636 3336 644 3344
rect 684 3336 692 3344
rect 956 3336 964 3344
rect 60 3318 68 3326
rect 124 3316 132 3324
rect 300 3318 308 3326
rect 1148 3336 1156 3344
rect 1180 3336 1188 3344
rect 1276 3336 1284 3344
rect 1612 3336 1620 3344
rect 1660 3336 1668 3344
rect 364 3316 372 3324
rect 476 3316 484 3324
rect 604 3316 612 3324
rect 636 3316 644 3324
rect 716 3316 724 3324
rect 764 3316 772 3324
rect 828 3316 836 3324
rect 908 3316 916 3324
rect 972 3316 980 3324
rect 1036 3316 1044 3324
rect 1068 3316 1076 3324
rect 1132 3316 1140 3324
rect 1164 3316 1172 3324
rect 1196 3316 1204 3324
rect 1276 3316 1284 3324
rect 1292 3316 1300 3324
rect 1388 3316 1396 3324
rect 1660 3316 1668 3324
rect 1724 3336 1732 3344
rect 1884 3336 1892 3344
rect 2108 3336 2116 3344
rect 2156 3336 2164 3344
rect 2188 3336 2196 3344
rect 2204 3336 2212 3344
rect 2348 3336 2356 3344
rect 2364 3336 2372 3344
rect 2428 3336 2436 3344
rect 2780 3356 2788 3364
rect 2876 3356 2884 3364
rect 3772 3356 3780 3364
rect 2476 3336 2484 3344
rect 1740 3316 1748 3324
rect 1756 3316 1764 3324
rect 1820 3316 1828 3324
rect 1884 3316 1892 3324
rect 1964 3316 1972 3324
rect 2060 3316 2068 3324
rect 2636 3336 2644 3344
rect 2300 3316 2308 3324
rect 2348 3316 2356 3324
rect 2412 3316 2420 3324
rect 2508 3316 2516 3324
rect 2556 3316 2564 3324
rect 2876 3336 2884 3344
rect 2940 3336 2948 3344
rect 3100 3336 3108 3344
rect 3180 3336 3188 3344
rect 3260 3336 3268 3344
rect 3500 3336 3508 3344
rect 3532 3336 3540 3344
rect 3548 3336 3556 3344
rect 3596 3336 3604 3344
rect 3628 3336 3636 3344
rect 3660 3336 3668 3344
rect 2700 3316 2708 3324
rect 2908 3316 2916 3324
rect 2956 3316 2964 3324
rect 3356 3316 3364 3324
rect 3388 3316 3396 3324
rect 3532 3316 3540 3324
rect 3548 3316 3556 3324
rect 3612 3316 3620 3324
rect 3644 3316 3652 3324
rect 492 3296 500 3304
rect 668 3296 676 3304
rect 716 3296 724 3304
rect 780 3296 788 3304
rect 844 3296 852 3304
rect 1052 3296 1060 3304
rect 1228 3296 1236 3304
rect 1388 3296 1396 3304
rect 1420 3296 1428 3304
rect 1500 3296 1508 3304
rect 1516 3296 1524 3304
rect 2028 3296 2036 3304
rect 2060 3296 2068 3304
rect 2092 3296 2100 3304
rect 2220 3296 2228 3304
rect 2252 3296 2260 3304
rect 2332 3296 2340 3304
rect 2476 3296 2484 3304
rect 2636 3296 2644 3304
rect 2700 3296 2708 3304
rect 2812 3296 2820 3304
rect 2844 3296 2852 3304
rect 2988 3296 2996 3304
rect 3208 3296 3216 3304
rect 3228 3296 3236 3304
rect 3276 3296 3284 3304
rect 3368 3296 3376 3304
rect 3388 3296 3396 3304
rect 3452 3296 3460 3304
rect 3676 3296 3684 3304
rect 3772 3336 3780 3344
rect 3740 3316 3748 3324
rect 3772 3316 3780 3324
rect 3804 3336 3812 3344
rect 4060 3336 4068 3344
rect 4092 3336 4100 3344
rect 4140 3336 4148 3344
rect 4188 3336 4196 3344
rect 4476 3356 4484 3364
rect 4748 3356 4756 3364
rect 4236 3336 4244 3344
rect 4332 3336 4340 3344
rect 5020 3356 5028 3364
rect 5628 3356 5636 3364
rect 5660 3356 5668 3364
rect 5740 3356 5748 3364
rect 4844 3336 4852 3344
rect 5084 3336 5092 3344
rect 5116 3336 5124 3344
rect 5180 3336 5188 3344
rect 5228 3336 5236 3344
rect 5244 3336 5252 3344
rect 5292 3336 5300 3344
rect 5388 3336 5396 3344
rect 5420 3336 5428 3344
rect 5436 3336 5444 3344
rect 5548 3336 5556 3344
rect 5612 3336 5620 3344
rect 5756 3336 5764 3344
rect 5836 3336 5844 3344
rect 5868 3356 5876 3364
rect 5996 3356 6004 3364
rect 5884 3336 5892 3344
rect 5964 3336 5972 3344
rect 6012 3336 6020 3344
rect 6060 3336 6068 3344
rect 6140 3336 6148 3344
rect 6252 3336 6260 3344
rect 3852 3316 3860 3324
rect 3964 3316 3972 3324
rect 4172 3316 4180 3324
rect 3724 3296 3732 3304
rect 4060 3296 4068 3304
rect 4108 3296 4116 3304
rect 4156 3296 4164 3304
rect 4268 3296 4276 3304
rect 4316 3316 4324 3324
rect 4428 3316 4436 3324
rect 4604 3316 4612 3324
rect 4620 3316 4628 3324
rect 4796 3316 4804 3324
rect 4316 3296 4324 3304
rect 4956 3316 4964 3324
rect 5004 3316 5012 3324
rect 4844 3296 4852 3304
rect 5116 3296 5124 3304
rect 5164 3316 5172 3324
rect 5196 3296 5204 3304
rect 5308 3316 5316 3324
rect 5372 3316 5380 3324
rect 5404 3316 5412 3324
rect 5436 3316 5444 3324
rect 5484 3316 5492 3324
rect 5532 3316 5540 3324
rect 5580 3316 5588 3324
rect 5596 3316 5604 3324
rect 5708 3316 5716 3324
rect 5340 3296 5348 3304
rect 5464 3296 5472 3304
rect 5500 3296 5508 3304
rect 5564 3296 5572 3304
rect 5740 3296 5748 3304
rect 5852 3316 5860 3324
rect 5900 3316 5908 3324
rect 5948 3316 5956 3324
rect 6028 3316 6036 3324
rect 6108 3316 6116 3324
rect 6140 3316 6148 3324
rect 6204 3316 6212 3324
rect 5804 3296 5812 3304
rect 5932 3296 5940 3304
rect 6060 3296 6068 3304
rect 6076 3296 6084 3304
rect 6220 3296 6228 3304
rect 460 3276 468 3284
rect 588 3276 596 3284
rect 748 3276 756 3284
rect 1084 3276 1092 3284
rect 1340 3276 1348 3284
rect 1372 3276 1380 3284
rect 3692 3276 3700 3284
rect 6108 3276 6116 3284
rect 220 3256 228 3264
rect 1356 3256 1364 3264
rect 1724 3256 1732 3264
rect 444 3236 452 3244
rect 524 3236 532 3244
rect 604 3236 612 3244
rect 764 3236 772 3244
rect 796 3236 804 3244
rect 1068 3236 1076 3244
rect 2460 3236 2468 3244
rect 2492 3236 2500 3244
rect 2732 3236 2740 3244
rect 2780 3236 2788 3244
rect 3036 3236 3044 3244
rect 3244 3236 3252 3244
rect 5900 3236 5908 3244
rect 5996 3236 6004 3244
rect 6092 3236 6100 3244
rect 6156 3236 6164 3244
rect 1577 3206 1585 3214
rect 1587 3206 1595 3214
rect 1597 3206 1605 3214
rect 1607 3206 1615 3214
rect 4665 3206 4673 3214
rect 4675 3206 4683 3214
rect 4685 3206 4693 3214
rect 4695 3206 4703 3214
rect 188 3176 196 3184
rect 348 3176 356 3184
rect 412 3176 420 3184
rect 1836 3176 1844 3184
rect 1932 3176 1940 3184
rect 2332 3176 2340 3184
rect 3084 3176 3092 3184
rect 3340 3176 3348 3184
rect 3388 3176 3396 3184
rect 3676 3176 3684 3184
rect 4236 3176 4244 3184
rect 4396 3176 4404 3184
rect 4508 3176 4516 3184
rect 4892 3176 4900 3184
rect 5836 3176 5844 3184
rect 780 3156 788 3164
rect 1244 3156 1252 3164
rect 1580 3156 1588 3164
rect 1612 3156 1620 3164
rect 5084 3156 5092 3164
rect 6092 3156 6100 3164
rect 364 3136 372 3144
rect 428 3136 436 3144
rect 460 3136 468 3144
rect 556 3136 564 3144
rect 716 3136 724 3144
rect 796 3136 804 3144
rect 988 3136 996 3144
rect 1100 3136 1108 3144
rect 1196 3136 1204 3144
rect 1260 3136 1268 3144
rect 1484 3136 1492 3144
rect 2652 3136 2660 3144
rect 2860 3136 2868 3144
rect 3068 3136 3076 3144
rect 3660 3136 3668 3144
rect 3788 3136 3796 3144
rect 3980 3136 3988 3144
rect 4124 3136 4132 3144
rect 4524 3136 4532 3144
rect 4796 3136 4804 3144
rect 5500 3136 5508 3144
rect 5596 3136 5604 3144
rect 5916 3136 5924 3144
rect 220 3116 228 3124
rect 332 3116 340 3124
rect 412 3116 420 3124
rect 492 3116 500 3124
rect 588 3116 596 3124
rect 652 3116 660 3124
rect 828 3116 836 3124
rect 876 3116 884 3124
rect 956 3116 964 3124
rect 1228 3116 1236 3124
rect 1516 3116 1524 3124
rect 1564 3116 1572 3124
rect 1644 3116 1652 3124
rect 92 3096 100 3104
rect 220 3096 228 3104
rect 252 3096 260 3104
rect 284 3096 292 3104
rect 316 3096 324 3104
rect 348 3096 356 3104
rect 412 3096 420 3104
rect 572 3096 580 3104
rect 620 3096 628 3104
rect 700 3096 708 3104
rect 764 3096 772 3104
rect 812 3096 820 3104
rect 972 3096 980 3104
rect 1148 3096 1156 3104
rect 1180 3096 1188 3104
rect 1196 3096 1204 3104
rect 1244 3096 1252 3104
rect 1356 3096 1364 3104
rect 76 3076 84 3084
rect 204 3076 212 3084
rect 268 3076 276 3084
rect 524 3076 532 3084
rect 604 3076 612 3084
rect 636 3076 644 3084
rect 716 3076 724 3084
rect 748 3076 756 3084
rect 844 3076 852 3084
rect 924 3080 932 3088
rect 1532 3096 1540 3104
rect 1564 3096 1572 3104
rect 1644 3096 1652 3104
rect 1692 3116 1700 3124
rect 1788 3116 1796 3124
rect 1804 3116 1812 3124
rect 1900 3116 1908 3124
rect 2076 3116 2084 3124
rect 2284 3116 2292 3124
rect 2300 3116 2308 3124
rect 2364 3116 2372 3124
rect 2428 3116 2436 3124
rect 2684 3116 2692 3124
rect 2700 3116 2708 3124
rect 2828 3116 2836 3124
rect 3132 3116 3140 3124
rect 1932 3096 1940 3104
rect 1964 3096 1972 3104
rect 2092 3096 2100 3104
rect 2204 3096 2212 3104
rect 940 3076 948 3084
rect 1020 3076 1028 3084
rect 1052 3076 1060 3084
rect 1084 3076 1092 3084
rect 1212 3076 1220 3084
rect 1308 3076 1316 3084
rect 1516 3076 1524 3084
rect 1532 3076 1540 3084
rect 1564 3076 1572 3084
rect 1628 3076 1636 3084
rect 1724 3076 1732 3084
rect 1740 3076 1748 3084
rect 1772 3076 1780 3084
rect 1852 3076 1860 3084
rect 1980 3076 1988 3084
rect 284 3056 292 3064
rect 684 3056 692 3064
rect 876 3056 884 3064
rect 1868 3056 1876 3064
rect 2028 3076 2036 3084
rect 2188 3076 2196 3084
rect 2348 3076 2356 3084
rect 2412 3096 2420 3104
rect 2524 3096 2532 3104
rect 2604 3096 2612 3104
rect 2668 3096 2676 3104
rect 2700 3096 2708 3104
rect 2732 3096 2740 3104
rect 2860 3096 2868 3104
rect 2940 3094 2948 3102
rect 3116 3096 3124 3104
rect 3372 3116 3380 3124
rect 3708 3116 3716 3124
rect 3820 3116 3828 3124
rect 3884 3116 3892 3124
rect 4108 3116 4116 3124
rect 4172 3116 4180 3124
rect 4192 3116 4200 3124
rect 4380 3116 4388 3124
rect 4428 3116 4436 3124
rect 3324 3096 3332 3104
rect 3532 3096 3540 3104
rect 3644 3096 3652 3104
rect 3804 3096 3812 3104
rect 3868 3096 3876 3104
rect 3932 3096 3940 3104
rect 2476 3076 2484 3084
rect 2540 3076 2548 3084
rect 2620 3076 2628 3084
rect 2764 3076 2772 3084
rect 2876 3076 2884 3084
rect 3132 3076 3140 3084
rect 3228 3076 3236 3084
rect 3436 3076 3444 3084
rect 3644 3076 3652 3084
rect 2140 3056 2148 3064
rect 2364 3056 2372 3064
rect 2812 3056 2820 3064
rect 3148 3056 3156 3064
rect 3308 3056 3316 3064
rect 3436 3056 3444 3064
rect 3708 3076 3716 3084
rect 3740 3076 3748 3084
rect 3852 3076 3860 3084
rect 3884 3076 3892 3084
rect 4076 3096 4084 3104
rect 4204 3096 4212 3104
rect 4300 3096 4308 3104
rect 4348 3096 4356 3104
rect 4668 3094 4676 3102
rect 4780 3096 4788 3104
rect 4844 3116 4852 3124
rect 5276 3116 5284 3124
rect 5420 3116 5428 3124
rect 5452 3116 5460 3124
rect 5804 3116 5812 3124
rect 5004 3096 5012 3104
rect 5212 3094 5220 3102
rect 5276 3096 5284 3104
rect 5324 3096 5332 3104
rect 5420 3096 5428 3104
rect 5452 3096 5460 3104
rect 5468 3096 5476 3104
rect 5548 3096 5556 3104
rect 5628 3096 5636 3104
rect 5708 3096 5716 3104
rect 5788 3096 5796 3104
rect 5836 3096 5844 3104
rect 5884 3116 5892 3124
rect 5948 3116 5956 3124
rect 5980 3116 5988 3124
rect 6156 3116 6164 3124
rect 6236 3116 6244 3124
rect 6284 3116 6292 3124
rect 5916 3096 5924 3104
rect 6156 3096 6164 3104
rect 6188 3096 6196 3104
rect 4220 3076 4228 3084
rect 4268 3076 4276 3084
rect 4332 3076 4340 3084
rect 4460 3076 4468 3084
rect 4700 3076 4708 3084
rect 4764 3076 4772 3084
rect 4876 3076 4884 3084
rect 5020 3076 5028 3084
rect 5196 3076 5204 3084
rect 5324 3076 5332 3084
rect 5468 3076 5476 3084
rect 5484 3076 5492 3084
rect 5532 3076 5540 3084
rect 5756 3076 5764 3084
rect 5932 3076 5940 3084
rect 5980 3076 5988 3084
rect 6028 3076 6036 3084
rect 6076 3076 6084 3084
rect 6204 3076 6212 3084
rect 6220 3076 6228 3084
rect 3772 3056 3780 3064
rect 3804 3056 3812 3064
rect 4284 3056 4292 3064
rect 4316 3056 4324 3064
rect 4412 3056 4420 3064
rect 4476 3056 4484 3064
rect 4524 3056 4532 3064
rect 5340 3056 5348 3064
rect 5372 3056 5380 3064
rect 5404 3056 5412 3064
rect 5564 3056 5572 3064
rect 5596 3056 5604 3064
rect 5676 3056 5684 3064
rect 5692 3056 5700 3064
rect 5724 3056 5732 3064
rect 5788 3056 5796 3064
rect 6108 3056 6116 3064
rect 6124 3056 6132 3064
rect 6156 3056 6164 3064
rect 492 3036 500 3044
rect 556 3036 564 3044
rect 668 3036 676 3044
rect 892 3036 900 3044
rect 1516 3036 1524 3044
rect 1612 3036 1620 3044
rect 2076 3036 2084 3044
rect 2156 3036 2164 3044
rect 2268 3036 2276 3044
rect 2524 3036 2532 3044
rect 2604 3036 2612 3044
rect 2796 3036 2804 3044
rect 3452 3036 3460 3044
rect 4108 3036 4116 3044
rect 4380 3036 4388 3044
rect 4428 3036 4436 3044
rect 4492 3036 4500 3044
rect 4892 3036 4900 3044
rect 5612 3036 5620 3044
rect 5660 3036 5668 3044
rect 5740 3036 5748 3044
rect 5948 3036 5956 3044
rect 6012 3036 6020 3044
rect 6044 3036 6052 3044
rect 3113 3006 3121 3014
rect 3123 3006 3131 3014
rect 3133 3006 3141 3014
rect 3143 3006 3151 3014
rect 60 2976 68 2984
rect 252 2976 260 2984
rect 348 2976 356 2984
rect 428 2976 436 2984
rect 1500 2976 1508 2984
rect 1836 2976 1844 2984
rect 1980 2976 1988 2984
rect 2572 2976 2580 2984
rect 2684 2976 2692 2984
rect 2748 2976 2756 2984
rect 2844 2976 2852 2984
rect 3004 2976 3012 2984
rect 3260 2976 3268 2984
rect 3404 2976 3412 2984
rect 3468 2976 3476 2984
rect 3580 2976 3588 2984
rect 3756 2976 3764 2984
rect 3932 2976 3940 2984
rect 4316 2976 4324 2984
rect 4508 2976 4516 2984
rect 4652 2976 4660 2984
rect 4972 2976 4980 2984
rect 5180 2976 5188 2984
rect 5260 2976 5268 2984
rect 5404 2976 5412 2984
rect 5676 2976 5684 2984
rect 5772 2976 5780 2984
rect 6268 2976 6276 2984
rect 540 2956 548 2964
rect 556 2956 564 2964
rect 604 2956 612 2964
rect 700 2956 708 2964
rect 780 2956 788 2964
rect 796 2956 804 2964
rect 12 2936 20 2944
rect 76 2936 84 2944
rect 140 2936 148 2944
rect 28 2916 36 2924
rect 60 2916 68 2924
rect 92 2916 100 2924
rect 124 2916 132 2924
rect 156 2916 164 2924
rect 188 2916 196 2924
rect 220 2936 228 2944
rect 332 2936 340 2944
rect 380 2936 388 2944
rect 652 2936 660 2944
rect 812 2936 820 2944
rect 828 2936 836 2944
rect 892 2936 900 2944
rect 972 2936 980 2944
rect 1084 2956 1092 2964
rect 1116 2956 1124 2964
rect 1308 2956 1316 2964
rect 1388 2956 1396 2964
rect 1676 2956 1684 2964
rect 1772 2956 1780 2964
rect 1916 2956 1924 2964
rect 1932 2956 1940 2964
rect 2236 2956 2244 2964
rect 2588 2956 2596 2964
rect 2732 2956 2740 2964
rect 2908 2956 2916 2964
rect 2940 2956 2948 2964
rect 2988 2956 2996 2964
rect 3388 2956 3396 2964
rect 3724 2956 3732 2964
rect 3868 2956 3876 2964
rect 4604 2956 4612 2964
rect 5340 2956 5348 2964
rect 5420 2956 5428 2964
rect 5436 2956 5444 2964
rect 5500 2956 5508 2964
rect 5564 2956 5572 2964
rect 5964 2956 5972 2964
rect 6076 2956 6084 2964
rect 6236 2956 6244 2964
rect 6252 2956 6260 2964
rect 1084 2936 1092 2944
rect 1148 2936 1156 2944
rect 1228 2936 1236 2944
rect 1340 2936 1348 2944
rect 1484 2936 1492 2944
rect 1660 2936 1668 2944
rect 1692 2936 1700 2944
rect 1788 2936 1796 2944
rect 1804 2936 1812 2944
rect 1852 2936 1860 2944
rect 1948 2936 1956 2944
rect 1996 2936 2004 2944
rect 2108 2936 2116 2944
rect 2236 2936 2244 2944
rect 2620 2936 2628 2944
rect 2636 2936 2644 2944
rect 2716 2936 2724 2944
rect 2764 2936 2772 2944
rect 2780 2936 2788 2944
rect 2796 2936 2804 2944
rect 3020 2936 3028 2944
rect 3228 2936 3236 2944
rect 3276 2936 3284 2944
rect 3308 2936 3316 2944
rect 3324 2936 3332 2944
rect 3356 2936 3364 2944
rect 3452 2936 3460 2944
rect 3532 2936 3540 2944
rect 3676 2936 3684 2944
rect 3804 2936 3812 2944
rect 3916 2936 3924 2944
rect 156 2896 164 2904
rect 300 2916 308 2924
rect 396 2916 404 2924
rect 460 2916 468 2924
rect 508 2916 516 2924
rect 604 2916 612 2924
rect 668 2916 676 2924
rect 748 2916 756 2924
rect 876 2916 884 2924
rect 940 2916 948 2924
rect 972 2916 980 2924
rect 1036 2916 1044 2924
rect 1068 2916 1076 2924
rect 1164 2916 1172 2924
rect 1180 2916 1188 2924
rect 1260 2916 1268 2924
rect 1356 2916 1364 2924
rect 1436 2916 1444 2924
rect 1532 2916 1540 2924
rect 1628 2916 1636 2924
rect 1788 2916 1796 2924
rect 2076 2916 2084 2924
rect 2108 2916 2116 2924
rect 2124 2916 2132 2924
rect 2268 2916 2276 2924
rect 2316 2916 2324 2924
rect 2380 2916 2388 2924
rect 2460 2916 2468 2924
rect 2812 2916 2820 2924
rect 2956 2916 2964 2924
rect 3164 2916 3172 2924
rect 3404 2916 3412 2924
rect 3436 2916 3444 2924
rect 3500 2916 3508 2924
rect 3596 2916 3604 2924
rect 3660 2916 3668 2924
rect 3820 2916 3828 2924
rect 3900 2916 3908 2924
rect 3948 2916 3956 2924
rect 3964 2916 3972 2924
rect 3980 2916 3988 2924
rect 4028 2916 4036 2924
rect 4172 2936 4180 2944
rect 4268 2936 4276 2944
rect 4284 2936 4292 2944
rect 4380 2936 4388 2944
rect 4524 2936 4532 2944
rect 4540 2936 4548 2944
rect 4556 2936 4564 2944
rect 5020 2936 5028 2944
rect 5164 2936 5172 2944
rect 5212 2936 5220 2944
rect 5276 2936 5284 2944
rect 5308 2936 5316 2944
rect 5388 2936 5396 2944
rect 5516 2936 5524 2944
rect 5628 2936 5636 2944
rect 5660 2936 5668 2944
rect 5692 2936 5700 2944
rect 5724 2936 5732 2944
rect 5980 2936 5988 2944
rect 6028 2936 6036 2944
rect 6044 2936 6052 2944
rect 6156 2936 6164 2944
rect 6220 2936 6228 2944
rect 4396 2916 4404 2924
rect 4572 2916 4580 2924
rect 4636 2916 4644 2924
rect 4732 2916 4740 2924
rect 4860 2916 4868 2924
rect 316 2896 324 2904
rect 364 2896 372 2904
rect 716 2896 724 2904
rect 736 2896 744 2904
rect 956 2896 964 2904
rect 988 2896 996 2904
rect 1100 2896 1108 2904
rect 1244 2896 1252 2904
rect 2044 2896 2052 2904
rect 2684 2896 2692 2904
rect 2860 2896 2868 2904
rect 2892 2896 2900 2904
rect 3052 2896 3060 2904
rect 3404 2896 3412 2904
rect 3468 2896 3476 2904
rect 3708 2896 3716 2904
rect 3852 2896 3860 2904
rect 4012 2896 4020 2904
rect 4316 2896 4324 2904
rect 4556 2896 4564 2904
rect 4620 2896 4628 2904
rect 5020 2896 5028 2904
rect 5068 2916 5076 2924
rect 5148 2916 5156 2924
rect 5212 2916 5220 2924
rect 5292 2916 5300 2924
rect 5516 2916 5524 2924
rect 5532 2916 5540 2924
rect 5116 2896 5124 2904
rect 5196 2896 5204 2904
rect 5260 2896 5268 2904
rect 5324 2896 5332 2904
rect 5612 2916 5620 2924
rect 5644 2916 5652 2924
rect 5708 2916 5716 2924
rect 5740 2916 5748 2924
rect 5804 2916 5812 2924
rect 5884 2916 5892 2924
rect 5980 2916 5988 2924
rect 6124 2916 6132 2924
rect 6172 2916 6180 2924
rect 5580 2896 5588 2904
rect 5772 2896 5780 2904
rect 5788 2896 5796 2904
rect 5900 2896 5908 2904
rect 6028 2896 6036 2904
rect 6076 2896 6084 2904
rect 6140 2896 6148 2904
rect 6204 2896 6212 2904
rect 220 2876 228 2884
rect 252 2876 260 2884
rect 284 2876 292 2884
rect 476 2876 484 2884
rect 924 2876 932 2884
rect 1276 2876 1284 2884
rect 1308 2876 1316 2884
rect 2188 2876 2196 2884
rect 2380 2876 2388 2884
rect 4092 2876 4100 2884
rect 4652 2876 4660 2884
rect 5468 2876 5476 2884
rect 5820 2876 5828 2884
rect 6108 2876 6116 2884
rect 908 2856 916 2864
rect 1628 2856 1636 2864
rect 492 2836 500 2844
rect 508 2836 516 2844
rect 668 2836 676 2844
rect 1116 2836 1124 2844
rect 1260 2836 1268 2844
rect 1500 2836 1508 2844
rect 2156 2836 2164 2844
rect 2268 2836 2276 2844
rect 2940 2836 2948 2844
rect 3084 2836 3092 2844
rect 3692 2836 3700 2844
rect 3836 2836 3844 2844
rect 4764 2836 4772 2844
rect 5804 2836 5812 2844
rect 5884 2836 5892 2844
rect 6124 2836 6132 2844
rect 6172 2836 6180 2844
rect 1577 2806 1585 2814
rect 1587 2806 1595 2814
rect 1597 2806 1605 2814
rect 1607 2806 1615 2814
rect 4665 2806 4673 2814
rect 4675 2806 4683 2814
rect 4685 2806 4693 2814
rect 4695 2806 4703 2814
rect 1100 2776 1108 2784
rect 1228 2776 1236 2784
rect 2012 2776 2020 2784
rect 2140 2776 2148 2784
rect 2428 2776 2436 2784
rect 2572 2776 2580 2784
rect 2876 2776 2884 2784
rect 2956 2776 2964 2784
rect 3164 2776 3172 2784
rect 3404 2776 3412 2784
rect 3516 2776 3524 2784
rect 3580 2776 3588 2784
rect 3660 2776 3668 2784
rect 3724 2776 3732 2784
rect 3900 2776 3908 2784
rect 4284 2776 4292 2784
rect 5468 2776 5476 2784
rect 5756 2776 5764 2784
rect 6012 2776 6020 2784
rect 6156 2776 6164 2784
rect 6204 2776 6212 2784
rect 220 2756 228 2764
rect 892 2756 900 2764
rect 956 2756 964 2764
rect 1324 2756 1332 2764
rect 3948 2756 3956 2764
rect 4076 2756 4084 2764
rect 252 2736 260 2744
rect 428 2736 436 2744
rect 444 2736 452 2744
rect 876 2736 884 2744
rect 940 2736 948 2744
rect 1084 2736 1092 2744
rect 1148 2736 1156 2744
rect 1212 2736 1220 2744
rect 1820 2736 1828 2744
rect 3004 2736 3012 2744
rect 3068 2736 3076 2744
rect 4044 2736 4052 2744
rect 5580 2736 5588 2744
rect 6140 2736 6148 2744
rect 188 2716 196 2724
rect 284 2716 292 2724
rect 556 2716 564 2724
rect 956 2716 964 2724
rect 1004 2716 1012 2724
rect 1116 2716 1124 2724
rect 1180 2716 1188 2724
rect 1244 2716 1252 2724
rect 1516 2716 1524 2724
rect 1596 2716 1604 2724
rect 2044 2716 2052 2724
rect 2108 2716 2116 2724
rect 2172 2716 2180 2724
rect 2220 2716 2228 2724
rect 2284 2716 2292 2724
rect 2332 2716 2340 2724
rect 2444 2716 2452 2724
rect 2508 2716 2516 2724
rect 2540 2716 2548 2724
rect 2924 2716 2932 2724
rect 3036 2716 3044 2724
rect 3100 2716 3108 2724
rect 3228 2716 3236 2724
rect 3324 2716 3332 2724
rect 3788 2716 3796 2724
rect 3852 2716 3860 2724
rect 4524 2716 4532 2724
rect 5148 2716 5156 2724
rect 5256 2716 5264 2724
rect 5276 2716 5284 2724
rect 76 2696 84 2704
rect 172 2696 180 2704
rect 220 2696 228 2704
rect 332 2696 340 2704
rect 348 2696 356 2704
rect 380 2696 388 2704
rect 412 2696 420 2704
rect 460 2696 468 2704
rect 572 2696 580 2704
rect 636 2696 644 2704
rect 668 2696 676 2704
rect 748 2694 756 2702
rect 956 2696 964 2704
rect 1052 2696 1060 2704
rect 1084 2696 1092 2704
rect 1132 2696 1140 2704
rect 1228 2696 1236 2704
rect 1308 2696 1316 2704
rect 1356 2696 1364 2704
rect 1388 2696 1396 2704
rect 1452 2696 1460 2704
rect 1548 2696 1556 2704
rect 1612 2696 1620 2704
rect 1644 2696 1652 2704
rect 1676 2696 1684 2704
rect 1772 2696 1780 2704
rect 1788 2696 1796 2704
rect 1916 2696 1924 2704
rect 1932 2696 1940 2704
rect 1996 2696 2004 2704
rect 2012 2696 2020 2704
rect 2124 2696 2132 2704
rect 92 2676 100 2684
rect 172 2676 180 2684
rect 236 2676 244 2684
rect 332 2676 340 2684
rect 364 2676 372 2684
rect 396 2676 404 2684
rect 492 2676 500 2684
rect 524 2676 532 2684
rect 652 2676 660 2684
rect 684 2676 692 2684
rect 716 2676 724 2684
rect 908 2676 916 2684
rect 1036 2676 1044 2684
rect 1132 2676 1140 2684
rect 1292 2676 1300 2684
rect 1372 2676 1380 2684
rect 1404 2676 1412 2684
rect 1468 2676 1476 2684
rect 1660 2676 1668 2684
rect 1692 2676 1700 2684
rect 1804 2676 1812 2684
rect 1900 2676 1908 2684
rect 1964 2676 1972 2684
rect 2124 2676 2132 2684
rect 2268 2676 2276 2684
rect 2492 2676 2500 2684
rect 2556 2696 2564 2704
rect 2652 2696 2660 2704
rect 2684 2696 2692 2704
rect 2764 2696 2772 2704
rect 2956 2696 2964 2704
rect 3148 2696 3156 2704
rect 3260 2696 3268 2704
rect 3276 2696 3284 2704
rect 2540 2676 2548 2684
rect 2556 2676 2564 2684
rect 2620 2676 2628 2684
rect 2684 2676 2692 2684
rect 2988 2676 2996 2684
rect 3116 2676 3124 2684
rect 3148 2676 3156 2684
rect 3276 2676 3284 2684
rect 140 2656 148 2664
rect 268 2656 276 2664
rect 604 2656 612 2664
rect 748 2656 756 2664
rect 1260 2656 1268 2664
rect 1436 2656 1444 2664
rect 1484 2656 1492 2664
rect 3324 2696 3332 2704
rect 3356 2696 3364 2704
rect 3404 2696 3412 2704
rect 3692 2696 3700 2704
rect 3756 2696 3764 2704
rect 3804 2696 3812 2704
rect 3820 2696 3828 2704
rect 4012 2696 4020 2704
rect 4268 2696 4276 2704
rect 4396 2696 4404 2704
rect 4492 2696 4500 2704
rect 4588 2694 4596 2702
rect 4652 2696 4660 2704
rect 4780 2696 4788 2704
rect 4796 2696 4804 2704
rect 4972 2696 4980 2704
rect 5020 2696 5028 2704
rect 5100 2696 5108 2704
rect 5116 2696 5124 2704
rect 5244 2696 5252 2704
rect 5340 2694 5348 2702
rect 5564 2696 5572 2704
rect 5628 2716 5636 2724
rect 5724 2716 5732 2724
rect 5896 2716 5904 2724
rect 5916 2716 5924 2724
rect 5980 2716 5988 2724
rect 6076 2716 6084 2724
rect 5756 2696 5764 2704
rect 5788 2696 5796 2704
rect 5852 2696 5860 2704
rect 5868 2696 5876 2704
rect 5932 2696 5940 2704
rect 6124 2696 6132 2704
rect 3372 2676 3380 2684
rect 3388 2676 3396 2684
rect 3452 2676 3460 2684
rect 3484 2676 3492 2684
rect 3532 2676 3540 2684
rect 3596 2676 3604 2684
rect 3612 2676 3620 2684
rect 3676 2676 3684 2684
rect 3836 2676 3844 2684
rect 3916 2676 3924 2684
rect 4012 2676 4020 2684
rect 4140 2676 4148 2684
rect 4236 2676 4244 2684
rect 4268 2676 4276 2684
rect 4380 2676 4388 2684
rect 4444 2676 4452 2684
rect 4476 2676 4484 2684
rect 4508 2676 4516 2684
rect 4844 2676 4852 2684
rect 5068 2676 5076 2684
rect 5228 2676 5236 2684
rect 5308 2676 5316 2684
rect 5548 2676 5556 2684
rect 5676 2676 5684 2684
rect 5772 2676 5780 2684
rect 5804 2676 5812 2684
rect 5852 2676 5860 2684
rect 5868 2676 5876 2684
rect 5932 2676 5940 2684
rect 6028 2676 6036 2684
rect 6108 2676 6116 2684
rect 6172 2716 6180 2724
rect 6236 2716 6244 2724
rect 6204 2696 6212 2704
rect 6188 2676 6196 2684
rect 3500 2656 3508 2664
rect 3868 2656 3876 2664
rect 3884 2656 3892 2664
rect 4892 2656 4900 2664
rect 5212 2656 5220 2664
rect 5484 2656 5492 2664
rect 5548 2656 5556 2664
rect 5692 2656 5700 2664
rect 5980 2656 5988 2664
rect 6044 2656 6052 2664
rect 6076 2656 6084 2664
rect 92 2636 100 2644
rect 284 2636 292 2644
rect 508 2636 516 2644
rect 556 2636 564 2644
rect 1276 2636 1284 2644
rect 1420 2636 1428 2644
rect 1708 2636 1716 2644
rect 2204 2636 2212 2644
rect 2364 2636 2372 2644
rect 2908 2636 2916 2644
rect 3036 2636 3044 2644
rect 3228 2636 3236 2644
rect 3324 2636 3332 2644
rect 3516 2636 3524 2644
rect 4172 2636 4180 2644
rect 4716 2636 4724 2644
rect 4908 2636 4916 2644
rect 5500 2636 5508 2644
rect 5708 2636 5716 2644
rect 5820 2636 5828 2644
rect 3113 2606 3121 2614
rect 3123 2606 3131 2614
rect 3133 2606 3141 2614
rect 3143 2606 3151 2614
rect 156 2576 164 2584
rect 540 2576 548 2584
rect 1292 2576 1300 2584
rect 2028 2576 2036 2584
rect 2092 2576 2100 2584
rect 2140 2576 2148 2584
rect 2172 2576 2180 2584
rect 2620 2576 2628 2584
rect 2684 2576 2692 2584
rect 3228 2576 3236 2584
rect 3356 2576 3364 2584
rect 3756 2576 3764 2584
rect 3884 2576 3892 2584
rect 4364 2576 4372 2584
rect 4764 2576 4772 2584
rect 5020 2576 5028 2584
rect 5484 2576 5492 2584
rect 6012 2576 6020 2584
rect 44 2556 52 2564
rect 76 2556 84 2564
rect 140 2556 148 2564
rect 252 2556 260 2564
rect 828 2556 836 2564
rect 1116 2556 1124 2564
rect 1228 2556 1236 2564
rect 1564 2556 1572 2564
rect 1916 2556 1924 2564
rect 2012 2556 2020 2564
rect 2156 2556 2164 2564
rect 2428 2556 2436 2564
rect 3004 2556 3012 2564
rect 3260 2556 3268 2564
rect 3372 2556 3380 2564
rect 3804 2556 3812 2564
rect 3932 2556 3940 2564
rect 4012 2556 4020 2564
rect 4652 2556 4660 2564
rect 5324 2556 5332 2564
rect 5340 2556 5348 2564
rect 92 2536 100 2544
rect 220 2536 228 2544
rect 332 2536 340 2544
rect 572 2536 580 2544
rect 636 2536 644 2544
rect 796 2536 804 2544
rect 876 2536 884 2544
rect 892 2536 900 2544
rect 940 2536 948 2544
rect 1148 2536 1156 2544
rect 1164 2536 1172 2544
rect 1324 2536 1332 2544
rect 1388 2536 1396 2544
rect 1548 2536 1556 2544
rect 1692 2536 1700 2544
rect 1724 2536 1732 2544
rect 1772 2536 1780 2544
rect 1868 2536 1876 2544
rect 2124 2536 2132 2544
rect 2412 2536 2420 2544
rect 2460 2536 2468 2544
rect 2572 2536 2580 2544
rect 2652 2536 2660 2544
rect 2700 2536 2708 2544
rect 2716 2536 2724 2544
rect 2780 2536 2788 2544
rect 2844 2536 2852 2544
rect 2860 2536 2868 2544
rect 2892 2536 2900 2544
rect 2924 2536 2932 2544
rect 2956 2536 2964 2544
rect 2988 2536 2996 2544
rect 3180 2536 3188 2544
rect 3244 2536 3252 2544
rect 3292 2536 3300 2544
rect 3308 2536 3316 2544
rect 12 2516 20 2524
rect 124 2516 132 2524
rect 188 2516 196 2524
rect 284 2516 292 2524
rect 300 2516 308 2524
rect 316 2516 324 2524
rect 396 2518 404 2526
rect 460 2516 468 2524
rect 540 2516 548 2524
rect 572 2516 580 2524
rect 620 2516 628 2524
rect 668 2516 676 2524
rect 716 2516 724 2524
rect 732 2516 740 2524
rect 748 2516 756 2524
rect 780 2516 788 2524
rect 844 2516 852 2524
rect 908 2516 916 2524
rect 972 2518 980 2526
rect 1148 2516 1156 2524
rect 1212 2516 1220 2524
rect 1260 2516 1268 2524
rect 1308 2516 1316 2524
rect 1372 2516 1380 2524
rect 1436 2516 1444 2524
rect 540 2496 548 2504
rect 588 2496 596 2504
rect 652 2496 660 2504
rect 764 2496 772 2504
rect 1196 2496 1204 2504
rect 1436 2496 1444 2504
rect 684 2476 692 2484
rect 1420 2476 1428 2484
rect 1484 2476 1492 2484
rect 1532 2516 1540 2524
rect 1676 2516 1684 2524
rect 1692 2516 1700 2524
rect 1788 2516 1796 2524
rect 1820 2516 1828 2524
rect 1884 2516 1892 2524
rect 2044 2516 2052 2524
rect 2108 2516 2116 2524
rect 2284 2516 2292 2524
rect 2396 2516 2404 2524
rect 2700 2516 2708 2524
rect 2732 2516 2740 2524
rect 2764 2516 2772 2524
rect 2796 2516 2804 2524
rect 2828 2516 2836 2524
rect 2876 2516 2884 2524
rect 2908 2516 2916 2524
rect 2940 2516 2948 2524
rect 3068 2516 3076 2524
rect 3196 2516 3204 2524
rect 3340 2536 3348 2544
rect 3580 2536 3588 2544
rect 3612 2536 3620 2544
rect 3644 2536 3652 2544
rect 3452 2516 3460 2524
rect 3788 2536 3796 2544
rect 3852 2536 3860 2544
rect 4044 2536 4052 2544
rect 4124 2536 4132 2544
rect 4332 2536 4340 2544
rect 4348 2536 4356 2544
rect 4444 2536 4452 2544
rect 4460 2536 4468 2544
rect 4572 2536 4580 2544
rect 4876 2536 4884 2544
rect 4988 2532 4996 2540
rect 5004 2536 5012 2544
rect 5276 2536 5284 2544
rect 5388 2536 5396 2544
rect 5996 2556 6004 2564
rect 5452 2536 5460 2544
rect 5484 2536 5492 2544
rect 5692 2536 5700 2544
rect 5724 2536 5732 2544
rect 5932 2536 5940 2544
rect 3852 2516 3860 2524
rect 3964 2516 3972 2524
rect 4012 2516 4020 2524
rect 4044 2516 4052 2524
rect 4060 2516 4068 2524
rect 4124 2516 4132 2524
rect 4204 2516 4212 2524
rect 4252 2516 4260 2524
rect 4268 2516 4276 2524
rect 4332 2516 4340 2524
rect 4428 2516 4436 2524
rect 4476 2516 4484 2524
rect 4524 2516 4532 2524
rect 4540 2516 4548 2524
rect 4636 2516 4644 2524
rect 4732 2516 4740 2524
rect 4748 2516 4756 2524
rect 4892 2518 4900 2526
rect 5084 2516 5092 2524
rect 5132 2516 5140 2524
rect 5212 2516 5220 2524
rect 5228 2516 5236 2524
rect 5420 2516 5428 2524
rect 5436 2516 5444 2524
rect 5500 2516 5508 2524
rect 5516 2516 5524 2524
rect 5628 2516 5636 2524
rect 5756 2516 5764 2524
rect 5916 2516 5924 2524
rect 6028 2516 6036 2524
rect 6156 2516 6164 2524
rect 6204 2516 6212 2524
rect 1516 2496 1524 2504
rect 1836 2496 1844 2504
rect 2092 2496 2100 2504
rect 3884 2496 3892 2504
rect 3916 2496 3924 2504
rect 3948 2496 3956 2504
rect 4076 2496 4084 2504
rect 4108 2496 4116 2504
rect 4140 2496 4148 2504
rect 4172 2496 4180 2504
rect 4284 2496 4292 2504
rect 4396 2496 4404 2504
rect 4508 2496 4516 2504
rect 4524 2496 4532 2504
rect 4956 2496 4964 2504
rect 5612 2496 5620 2504
rect 5708 2496 5716 2504
rect 5724 2496 5732 2504
rect 5788 2496 5796 2504
rect 6076 2496 6084 2504
rect 1516 2476 1524 2484
rect 2012 2476 2020 2484
rect 2396 2476 2404 2484
rect 3084 2476 3092 2484
rect 3116 2476 3124 2484
rect 3564 2476 3572 2484
rect 3980 2476 3988 2484
rect 5756 2476 5764 2484
rect 5804 2476 5812 2484
rect 6044 2476 6052 2484
rect 1132 2456 1140 2464
rect 1340 2456 1348 2464
rect 2828 2456 2836 2464
rect 1404 2436 1412 2444
rect 1500 2436 1508 2444
rect 1724 2436 1732 2444
rect 1820 2436 1828 2444
rect 1852 2436 1860 2444
rect 2444 2436 2452 2444
rect 3660 2436 3668 2444
rect 3836 2436 3844 2444
rect 3964 2436 3972 2444
rect 4300 2436 4308 2444
rect 5548 2436 5556 2444
rect 5596 2436 5604 2444
rect 6092 2436 6100 2444
rect 1577 2406 1585 2414
rect 1587 2406 1595 2414
rect 1597 2406 1605 2414
rect 1607 2406 1615 2414
rect 4665 2406 4673 2414
rect 4675 2406 4683 2414
rect 4685 2406 4693 2414
rect 4695 2406 4703 2414
rect 44 2376 52 2384
rect 844 2376 852 2384
rect 1372 2376 1380 2384
rect 1420 2376 1428 2384
rect 2524 2376 2532 2384
rect 2844 2376 2852 2384
rect 2988 2376 2996 2384
rect 3388 2376 3396 2384
rect 3564 2376 3572 2384
rect 4268 2376 4276 2384
rect 4316 2376 4324 2384
rect 4428 2376 4436 2384
rect 4508 2376 4516 2384
rect 5260 2376 5268 2384
rect 1308 2356 1316 2364
rect 860 2336 868 2344
rect 1244 2336 1252 2344
rect 1484 2336 1492 2344
rect 1724 2356 1732 2364
rect 2636 2356 2644 2364
rect 1516 2336 1524 2344
rect 1932 2336 1940 2344
rect 2876 2336 2884 2344
rect 3820 2336 3828 2344
rect 4124 2336 4132 2344
rect 4156 2336 4164 2344
rect 4380 2336 4388 2344
rect 4444 2336 4452 2344
rect 428 2316 436 2324
rect 524 2316 532 2324
rect 636 2316 644 2324
rect 716 2316 724 2324
rect 828 2316 836 2324
rect 1036 2316 1044 2324
rect 1276 2316 1284 2324
rect 1340 2316 1348 2324
rect 1452 2316 1460 2324
rect 1516 2316 1524 2324
rect 1788 2316 1796 2324
rect 1900 2316 1908 2324
rect 2172 2316 2180 2324
rect 2204 2316 2212 2324
rect 2220 2316 2228 2324
rect 2332 2316 2340 2324
rect 2780 2316 2788 2324
rect 2956 2316 2964 2324
rect 3596 2316 3604 2324
rect 12 2296 20 2304
rect 140 2296 148 2304
rect 188 2296 196 2304
rect 348 2296 356 2304
rect 380 2296 388 2304
rect 476 2296 484 2304
rect 556 2296 564 2304
rect 636 2296 644 2304
rect 732 2296 740 2304
rect 780 2296 788 2304
rect 812 2296 820 2304
rect 844 2296 852 2304
rect 892 2296 900 2304
rect 956 2296 964 2304
rect 972 2296 980 2304
rect 988 2296 996 2304
rect 1116 2296 1124 2304
rect 1324 2296 1332 2304
rect 1388 2296 1396 2304
rect 1500 2296 1508 2304
rect 1692 2296 1700 2304
rect 1788 2296 1796 2304
rect 1852 2296 1860 2304
rect 2092 2294 2100 2302
rect 2172 2296 2180 2304
rect 2412 2296 2420 2304
rect 2748 2296 2756 2304
rect 2876 2296 2884 2304
rect 2988 2296 2996 2304
rect 3292 2296 3300 2304
rect 3324 2296 3332 2304
rect 3356 2296 3364 2304
rect 3372 2296 3380 2304
rect 3564 2296 3572 2304
rect 3612 2296 3620 2304
rect 3676 2296 3684 2304
rect 4188 2316 4196 2324
rect 4348 2316 4356 2324
rect 4412 2316 4420 2324
rect 4524 2336 4532 2344
rect 5212 2336 5220 2344
rect 5244 2336 5252 2344
rect 6252 2336 6260 2344
rect 4492 2316 4500 2324
rect 5644 2316 5652 2324
rect 5740 2316 5748 2324
rect 3820 2296 3828 2304
rect 3868 2296 3876 2304
rect 3916 2296 3924 2304
rect 3932 2296 3940 2304
rect 3996 2294 4004 2302
rect 4156 2296 4164 2304
rect 4204 2296 4212 2304
rect 60 2276 68 2284
rect 268 2276 276 2284
rect 300 2276 308 2284
rect 332 2276 340 2284
rect 572 2276 580 2284
rect 668 2276 676 2284
rect 684 2276 692 2284
rect 748 2276 756 2284
rect 412 2256 420 2264
rect 428 2256 436 2264
rect 508 2256 516 2264
rect 620 2256 628 2264
rect 796 2276 804 2284
rect 940 2276 948 2284
rect 1068 2276 1076 2284
rect 1324 2276 1332 2284
rect 1388 2276 1396 2284
rect 1548 2276 1556 2284
rect 1580 2276 1588 2284
rect 1676 2276 1684 2284
rect 1708 2276 1716 2284
rect 1756 2276 1764 2284
rect 1820 2276 1828 2284
rect 2156 2276 2164 2284
rect 2268 2276 2276 2284
rect 2316 2276 2324 2284
rect 2556 2276 2564 2284
rect 2652 2276 2660 2284
rect 2716 2276 2724 2284
rect 2732 2276 2740 2284
rect 2796 2276 2804 2284
rect 3004 2276 3012 2284
rect 3260 2276 3268 2284
rect 3340 2276 3348 2284
rect 3372 2276 3380 2284
rect 3420 2276 3428 2284
rect 3516 2280 3524 2288
rect 3532 2276 3540 2284
rect 3548 2276 3556 2284
rect 3628 2276 3636 2284
rect 3692 2276 3700 2284
rect 3740 2276 3748 2284
rect 3852 2276 3860 2284
rect 4140 2276 4148 2284
rect 4236 2276 4244 2284
rect 4284 2276 4292 2284
rect 4316 2296 4324 2304
rect 4380 2296 4388 2304
rect 4444 2296 4452 2304
rect 4508 2296 4516 2304
rect 4668 2296 4676 2304
rect 4924 2296 4932 2304
rect 5116 2296 5124 2304
rect 5372 2296 5380 2304
rect 5516 2296 5524 2304
rect 5580 2294 5588 2302
rect 5644 2296 5652 2304
rect 5676 2296 5684 2304
rect 5820 2296 5828 2304
rect 6284 2316 6292 2324
rect 6108 2296 6116 2304
rect 6156 2296 6164 2304
rect 6252 2296 6260 2304
rect 4364 2276 4372 2284
rect 4716 2276 4724 2284
rect 4892 2276 4900 2284
rect 5084 2276 5092 2284
rect 5212 2276 5220 2284
rect 5420 2276 5428 2284
rect 5692 2276 5700 2284
rect 5708 2276 5716 2284
rect 5804 2276 5812 2284
rect 5820 2276 5828 2284
rect 5916 2276 5924 2284
rect 5932 2276 5940 2284
rect 5996 2276 6004 2284
rect 6028 2276 6036 2284
rect 796 2256 804 2264
rect 892 2256 900 2264
rect 924 2256 932 2264
rect 1020 2256 1028 2264
rect 1244 2256 1252 2264
rect 1724 2256 1732 2264
rect 1788 2256 1796 2264
rect 1852 2256 1860 2264
rect 2588 2256 2596 2264
rect 2668 2256 2676 2264
rect 2924 2256 2932 2264
rect 3308 2256 3316 2264
rect 3468 2256 3476 2264
rect 3644 2256 3652 2264
rect 3660 2256 3668 2264
rect 3724 2256 3732 2264
rect 4252 2256 4260 2264
rect 4796 2256 4804 2264
rect 4812 2256 4820 2264
rect 252 2236 260 2244
rect 524 2236 532 2244
rect 700 2236 708 2244
rect 1580 2236 1588 2244
rect 1964 2236 1972 2244
rect 2940 2236 2948 2244
rect 3020 2236 3028 2244
rect 3484 2236 3492 2244
rect 3708 2236 3716 2244
rect 4556 2236 4564 2244
rect 4828 2236 4836 2244
rect 5228 2236 5236 2244
rect 5260 2236 5268 2244
rect 5756 2236 5764 2244
rect 5852 2236 5860 2244
rect 6044 2236 6052 2244
rect 3113 2206 3121 2214
rect 3123 2206 3131 2214
rect 3133 2206 3141 2214
rect 3143 2206 3151 2214
rect 396 2176 404 2184
rect 684 2176 692 2184
rect 1084 2176 1092 2184
rect 1196 2176 1204 2184
rect 1948 2176 1956 2184
rect 2396 2176 2404 2184
rect 2412 2176 2420 2184
rect 2556 2176 2564 2184
rect 2748 2176 2756 2184
rect 2860 2176 2868 2184
rect 2892 2176 2900 2184
rect 3052 2176 3060 2184
rect 3212 2176 3220 2184
rect 3612 2176 3620 2184
rect 3692 2176 3700 2184
rect 4620 2176 4628 2184
rect 4780 2176 4788 2184
rect 4924 2176 4932 2184
rect 5020 2176 5028 2184
rect 5164 2176 5172 2184
rect 6012 2176 6020 2184
rect 6092 2176 6100 2184
rect 204 2156 212 2164
rect 812 2156 820 2164
rect 1020 2156 1028 2164
rect 1260 2156 1268 2164
rect 1404 2156 1412 2164
rect 1452 2156 1460 2164
rect 1708 2156 1716 2164
rect 1740 2156 1748 2164
rect 2156 2156 2164 2164
rect 2236 2156 2244 2164
rect 2476 2156 2484 2164
rect 2572 2156 2580 2164
rect 2652 2156 2660 2164
rect 2764 2156 2772 2164
rect 124 2136 132 2144
rect 252 2136 260 2144
rect 380 2136 388 2144
rect 428 2136 436 2144
rect 524 2136 532 2144
rect 700 2136 708 2144
rect 796 2136 804 2144
rect 908 2136 916 2144
rect 140 2118 148 2126
rect 268 2116 276 2124
rect 300 2116 308 2124
rect 364 2116 372 2124
rect 428 2116 436 2124
rect 460 2116 468 2124
rect 572 2116 580 2124
rect 716 2116 724 2124
rect 204 2096 212 2104
rect 316 2096 324 2104
rect 348 2096 356 2104
rect 716 2096 724 2104
rect 844 2116 852 2124
rect 860 2116 868 2124
rect 924 2116 932 2124
rect 972 2116 980 2124
rect 3484 2156 3492 2164
rect 1116 2136 1124 2144
rect 1244 2136 1252 2144
rect 1356 2136 1364 2144
rect 1372 2136 1380 2144
rect 1564 2136 1572 2144
rect 1580 2136 1588 2144
rect 1804 2136 1812 2144
rect 1884 2136 1892 2144
rect 2140 2136 2148 2144
rect 2188 2136 2196 2144
rect 2220 2136 2228 2144
rect 2348 2136 2356 2144
rect 2492 2136 2500 2144
rect 2604 2136 2612 2144
rect 2636 2136 2644 2144
rect 2700 2136 2708 2144
rect 2732 2136 2740 2144
rect 1068 2116 1076 2124
rect 1132 2116 1140 2124
rect 1180 2116 1188 2124
rect 1340 2116 1348 2124
rect 1388 2116 1396 2124
rect 1500 2116 1508 2124
rect 1676 2116 1684 2124
rect 1788 2116 1796 2124
rect 1820 2116 1828 2124
rect 2028 2116 2036 2124
rect 2044 2116 2052 2124
rect 2236 2116 2244 2124
rect 2268 2116 2276 2124
rect 2316 2116 2324 2124
rect 2364 2116 2372 2124
rect 2460 2116 2468 2124
rect 2652 2116 2660 2124
rect 2684 2116 2692 2124
rect 2812 2136 2820 2144
rect 2876 2136 2884 2144
rect 2940 2136 2948 2144
rect 3004 2136 3012 2144
rect 3116 2136 3124 2144
rect 3228 2136 3236 2144
rect 3468 2136 3476 2144
rect 3500 2136 3508 2144
rect 3516 2136 3524 2144
rect 3756 2156 3764 2164
rect 3820 2156 3828 2164
rect 4204 2156 4212 2164
rect 4268 2156 4276 2164
rect 4588 2156 4596 2164
rect 4700 2156 4708 2164
rect 4796 2156 4804 2164
rect 5004 2156 5012 2164
rect 5180 2156 5188 2164
rect 5516 2156 5524 2164
rect 5676 2156 5684 2164
rect 3628 2136 3636 2144
rect 3788 2136 3796 2144
rect 3852 2136 3860 2144
rect 3868 2136 3876 2144
rect 3932 2136 3940 2144
rect 3948 2136 3956 2144
rect 4204 2136 4212 2144
rect 4236 2136 4244 2144
rect 4300 2136 4308 2144
rect 4444 2136 4452 2144
rect 4588 2136 4596 2144
rect 4716 2136 4724 2144
rect 4732 2136 4740 2144
rect 4860 2136 4868 2144
rect 4876 2136 4884 2144
rect 4988 2136 4996 2144
rect 5052 2136 5060 2144
rect 5084 2136 5092 2144
rect 5116 2136 5124 2144
rect 5356 2136 5364 2144
rect 5500 2136 5508 2144
rect 5596 2136 5604 2144
rect 2812 2116 2820 2124
rect 2860 2116 2868 2124
rect 2940 2116 2948 2124
rect 2988 2116 2996 2124
rect 3020 2116 3028 2124
rect 3036 2116 3044 2124
rect 3164 2116 3172 2124
rect 3180 2116 3188 2124
rect 3372 2116 3380 2124
rect 3452 2116 3460 2124
rect 3532 2116 3540 2124
rect 3580 2116 3588 2124
rect 3644 2116 3652 2124
rect 3692 2116 3700 2124
rect 3724 2116 3732 2124
rect 3804 2116 3812 2124
rect 764 2096 772 2104
rect 972 2096 980 2104
rect 476 2076 484 2084
rect 956 2076 964 2084
rect 1196 2096 1204 2104
rect 1452 2096 1460 2104
rect 1516 2096 1524 2104
rect 1644 2096 1652 2104
rect 1996 2096 2004 2104
rect 2108 2096 2116 2104
rect 2332 2096 2340 2104
rect 2588 2096 2596 2104
rect 2652 2096 2660 2104
rect 2780 2096 2788 2104
rect 2892 2096 2900 2104
rect 2956 2096 2964 2104
rect 3212 2096 3220 2104
rect 3612 2096 3620 2104
rect 3676 2096 3684 2104
rect 3692 2096 3700 2104
rect 3884 2116 3892 2124
rect 3916 2116 3924 2124
rect 3964 2116 3972 2124
rect 3980 2116 3988 2124
rect 4060 2118 4068 2126
rect 4252 2116 4260 2124
rect 4364 2116 4372 2124
rect 4412 2116 4420 2124
rect 4428 2116 4436 2124
rect 4460 2116 4468 2124
rect 4556 2116 4564 2124
rect 4748 2116 4756 2124
rect 3916 2096 3924 2104
rect 3996 2096 4004 2104
rect 4284 2096 4292 2104
rect 4332 2096 4340 2104
rect 4380 2096 4388 2104
rect 4472 2096 4480 2104
rect 4828 2116 4836 2124
rect 4876 2116 4884 2124
rect 4924 2116 4932 2124
rect 5036 2116 5044 2124
rect 5068 2116 5076 2124
rect 5324 2118 5332 2126
rect 5468 2116 5476 2124
rect 5676 2116 5684 2124
rect 5740 2118 5748 2126
rect 5804 2116 5812 2124
rect 5852 2116 5860 2124
rect 6076 2136 6084 2144
rect 6012 2116 6020 2124
rect 6156 2116 6164 2124
rect 6204 2116 6212 2124
rect 5148 2096 5156 2104
rect 492 2056 500 2064
rect 1036 2076 1044 2084
rect 1148 2076 1156 2084
rect 2172 2076 2180 2084
rect 5836 2076 5844 2084
rect 5916 2076 5924 2084
rect 5388 2056 5396 2064
rect 828 2036 836 2044
rect 876 2036 884 2044
rect 1020 2036 1028 2044
rect 1468 2036 1476 2044
rect 1836 2036 1844 2044
rect 3260 2036 3268 2044
rect 3548 2036 3556 2044
rect 4188 2036 4196 2044
rect 4844 2036 4852 2044
rect 5196 2036 5204 2044
rect 5580 2036 5588 2044
rect 5612 2036 5620 2044
rect 1577 2006 1585 2014
rect 1587 2006 1595 2014
rect 1597 2006 1605 2014
rect 1607 2006 1615 2014
rect 4665 2006 4673 2014
rect 4675 2006 4683 2014
rect 4685 2006 4693 2014
rect 4695 2006 4703 2014
rect 12 1976 20 1984
rect 492 1976 500 1984
rect 636 1976 644 1984
rect 1148 1976 1156 1984
rect 1356 1976 1364 1984
rect 1660 1976 1668 1984
rect 1692 1976 1700 1984
rect 1772 1976 1780 1984
rect 2044 1976 2052 1984
rect 2300 1976 2308 1984
rect 2396 1976 2404 1984
rect 2572 1976 2580 1984
rect 2620 1976 2628 1984
rect 3020 1976 3028 1984
rect 3068 1976 3076 1984
rect 3452 1976 3460 1984
rect 3692 1976 3700 1984
rect 3788 1976 3796 1984
rect 3836 1976 3844 1984
rect 3948 1976 3956 1984
rect 4028 1976 4036 1984
rect 4652 1976 4660 1984
rect 4908 1976 4916 1984
rect 4988 1976 4996 1984
rect 5036 1976 5044 1984
rect 6060 1976 6068 1984
rect 6188 1976 6196 1984
rect 428 1956 436 1964
rect 1068 1956 1076 1964
rect 2412 1956 2420 1964
rect 4348 1956 4356 1964
rect 5164 1956 5172 1964
rect 5932 1956 5940 1964
rect 6156 1956 6164 1964
rect 444 1936 452 1944
rect 572 1936 580 1944
rect 1276 1936 1284 1944
rect 1996 1936 2004 1944
rect 2236 1936 2244 1944
rect 2316 1936 2324 1944
rect 2716 1936 2724 1944
rect 2940 1936 2948 1944
rect 3724 1936 3732 1944
rect 4252 1936 4260 1944
rect 4300 1936 4308 1944
rect 4636 1936 4644 1944
rect 5212 1936 5220 1944
rect 5244 1936 5252 1944
rect 5324 1936 5332 1944
rect 5500 1936 5508 1944
rect 6108 1936 6116 1944
rect 6204 1936 6212 1944
rect 284 1916 292 1924
rect 396 1916 404 1924
rect 412 1916 420 1924
rect 540 1916 548 1924
rect 652 1916 660 1924
rect 716 1916 724 1924
rect 736 1916 744 1924
rect 972 1916 980 1924
rect 1180 1916 1188 1924
rect 1516 1916 1524 1924
rect 1980 1916 1988 1924
rect 2140 1916 2148 1924
rect 2348 1916 2356 1924
rect 2684 1916 2692 1924
rect 2796 1916 2804 1924
rect 3276 1916 3284 1924
rect 3324 1916 3332 1924
rect 3388 1916 3396 1924
rect 3516 1916 3524 1924
rect 3580 1916 3588 1924
rect 3740 1916 3748 1924
rect 3756 1916 3764 1924
rect 3868 1916 3876 1924
rect 3964 1916 3972 1924
rect 4092 1916 4100 1924
rect 4108 1916 4116 1924
rect 4128 1916 4136 1924
rect 4188 1916 4196 1924
rect 4220 1916 4228 1924
rect 4604 1916 4612 1924
rect 4828 1916 4836 1924
rect 4940 1916 4948 1924
rect 4956 1916 4964 1924
rect 5068 1916 5076 1924
rect 5084 1916 5092 1924
rect 5196 1916 5204 1924
rect 5340 1916 5348 1924
rect 5360 1916 5368 1924
rect 5404 1916 5412 1924
rect 6028 1916 6036 1924
rect 6140 1916 6148 1924
rect 140 1894 148 1902
rect 204 1896 212 1904
rect 284 1896 292 1904
rect 348 1896 356 1904
rect 364 1896 372 1904
rect 428 1896 436 1904
rect 588 1896 596 1904
rect 604 1896 612 1904
rect 684 1896 692 1904
rect 748 1896 756 1904
rect 844 1896 852 1904
rect 1020 1896 1028 1904
rect 1132 1896 1140 1904
rect 1228 1896 1236 1904
rect 1276 1896 1284 1904
rect 1324 1896 1332 1904
rect 1372 1896 1380 1904
rect 1452 1896 1460 1904
rect 1644 1896 1652 1904
rect 124 1876 132 1884
rect 172 1876 180 1884
rect 220 1876 228 1884
rect 332 1876 340 1884
rect 348 1876 356 1884
rect 476 1876 484 1884
rect 508 1876 516 1884
rect 668 1876 676 1884
rect 700 1876 708 1884
rect 764 1876 772 1884
rect 796 1876 804 1884
rect 972 1876 980 1884
rect 1100 1876 1108 1884
rect 1132 1876 1140 1884
rect 1244 1876 1252 1884
rect 1260 1876 1268 1884
rect 1324 1876 1332 1884
rect 1388 1876 1396 1884
rect 1436 1876 1444 1884
rect 1468 1876 1476 1884
rect 1548 1876 1556 1884
rect 1612 1876 1620 1884
rect 1900 1896 1908 1904
rect 1948 1896 1956 1904
rect 1980 1896 1988 1904
rect 2044 1896 2052 1904
rect 2156 1896 2164 1904
rect 252 1856 260 1864
rect 620 1856 628 1864
rect 1052 1856 1060 1864
rect 1068 1856 1076 1864
rect 1404 1856 1412 1864
rect 1532 1856 1540 1864
rect 1692 1856 1700 1864
rect 1804 1856 1812 1864
rect 1916 1876 1924 1884
rect 2028 1876 2036 1884
rect 2156 1876 2164 1884
rect 1916 1856 1924 1864
rect 1980 1856 1988 1864
rect 2156 1856 2164 1864
rect 2236 1896 2244 1904
rect 2252 1896 2260 1904
rect 2332 1896 2340 1904
rect 2396 1896 2404 1904
rect 2460 1896 2468 1904
rect 2636 1896 2644 1904
rect 2700 1896 2708 1904
rect 2780 1896 2788 1904
rect 2812 1896 2820 1904
rect 2988 1896 2996 1904
rect 3036 1896 3044 1904
rect 3180 1896 3188 1904
rect 3196 1896 3204 1904
rect 3388 1896 3396 1904
rect 3404 1896 3412 1904
rect 3548 1896 3556 1904
rect 3676 1896 3684 1904
rect 3724 1896 3732 1904
rect 3772 1896 3780 1904
rect 3804 1896 3812 1904
rect 3836 1896 3844 1904
rect 3868 1896 3876 1904
rect 3932 1896 3940 1904
rect 3980 1896 3988 1904
rect 4044 1896 4052 1904
rect 4108 1896 4116 1904
rect 4140 1896 4148 1904
rect 4188 1896 4196 1904
rect 4252 1896 4260 1904
rect 4460 1896 4468 1904
rect 4540 1896 4548 1904
rect 4684 1896 4692 1904
rect 4764 1896 4772 1904
rect 4780 1896 4788 1904
rect 4812 1896 4820 1904
rect 4860 1896 4868 1904
rect 4892 1896 4900 1904
rect 4908 1896 4916 1904
rect 4988 1896 4996 1904
rect 5036 1896 5044 1904
rect 5116 1896 5124 1904
rect 5132 1896 5140 1904
rect 5244 1896 5252 1904
rect 5372 1896 5380 1904
rect 5420 1896 5428 1904
rect 5436 1896 5444 1904
rect 5548 1896 5556 1904
rect 5708 1896 5716 1904
rect 5820 1896 5828 1904
rect 5980 1896 5988 1904
rect 5996 1896 6004 1904
rect 6060 1896 6068 1904
rect 2284 1876 2292 1884
rect 2508 1876 2516 1884
rect 2892 1876 2900 1884
rect 2956 1876 2964 1884
rect 3148 1876 3156 1884
rect 3212 1876 3220 1884
rect 3292 1876 3300 1884
rect 3340 1876 3348 1884
rect 3436 1876 3444 1884
rect 2204 1856 2212 1864
rect 2284 1856 2292 1864
rect 2364 1856 2372 1864
rect 2476 1856 2484 1864
rect 2604 1856 2612 1864
rect 2812 1856 2820 1864
rect 3404 1856 3412 1864
rect 3436 1856 3444 1864
rect 3564 1876 3572 1884
rect 3612 1876 3620 1884
rect 3804 1876 3812 1884
rect 3820 1876 3828 1884
rect 3932 1876 3940 1884
rect 3996 1876 4004 1884
rect 4044 1876 4052 1884
rect 4156 1876 4164 1884
rect 4236 1876 4244 1884
rect 4332 1876 4340 1884
rect 4556 1876 4564 1884
rect 4732 1876 4740 1884
rect 4764 1876 4772 1884
rect 4876 1876 4884 1884
rect 5004 1876 5012 1884
rect 5020 1876 5028 1884
rect 5132 1876 5140 1884
rect 5148 1876 5156 1884
rect 5260 1876 5268 1884
rect 5324 1876 5332 1884
rect 5388 1876 5396 1884
rect 5452 1876 5460 1884
rect 5532 1876 5540 1884
rect 5676 1876 5684 1884
rect 5772 1876 5780 1884
rect 6076 1876 6084 1884
rect 6092 1876 6100 1884
rect 6252 1876 6260 1884
rect 4028 1856 4036 1864
rect 4588 1856 4596 1864
rect 4764 1856 4772 1864
rect 4812 1856 4820 1864
rect 5084 1856 5092 1864
rect 5740 1856 5748 1864
rect 5948 1856 5956 1864
rect 6012 1856 6020 1864
rect 6028 1856 6036 1864
rect 6172 1856 6180 1864
rect 6204 1856 6212 1864
rect 6268 1856 6276 1864
rect 396 1836 404 1844
rect 540 1836 548 1844
rect 588 1836 596 1844
rect 956 1836 964 1844
rect 1196 1836 1204 1844
rect 1420 1836 1428 1844
rect 1516 1836 1524 1844
rect 2572 1836 2580 1844
rect 2652 1836 2660 1844
rect 2764 1836 2772 1844
rect 3596 1836 3604 1844
rect 4300 1836 4308 1844
rect 4572 1836 4580 1844
rect 5468 1836 5476 1844
rect 5724 1836 5732 1844
rect 3113 1806 3121 1814
rect 3123 1806 3131 1814
rect 3133 1806 3141 1814
rect 3143 1806 3151 1814
rect 76 1776 84 1784
rect 220 1776 228 1784
rect 428 1776 436 1784
rect 620 1776 628 1784
rect 684 1776 692 1784
rect 988 1776 996 1784
rect 1068 1776 1076 1784
rect 1436 1776 1444 1784
rect 1628 1776 1636 1784
rect 1980 1776 1988 1784
rect 2012 1776 2020 1784
rect 2188 1776 2196 1784
rect 2396 1776 2404 1784
rect 2972 1776 2980 1784
rect 2988 1776 2996 1784
rect 3276 1776 3284 1784
rect 3324 1776 3332 1784
rect 3388 1776 3396 1784
rect 3756 1776 3764 1784
rect 4092 1776 4100 1784
rect 4124 1776 4132 1784
rect 4892 1776 4900 1784
rect 4940 1776 4948 1784
rect 5004 1776 5012 1784
rect 5052 1776 5060 1784
rect 5116 1776 5124 1784
rect 5612 1776 5620 1784
rect 5660 1776 5668 1784
rect 6076 1776 6084 1784
rect 60 1756 68 1764
rect 556 1756 564 1764
rect 780 1756 788 1764
rect 796 1756 804 1764
rect 828 1756 836 1764
rect 940 1756 948 1764
rect 1484 1756 1492 1764
rect 1612 1756 1620 1764
rect 1676 1756 1684 1764
rect 28 1736 36 1744
rect 124 1736 132 1744
rect 236 1736 244 1744
rect 2028 1756 2036 1764
rect 2204 1756 2212 1764
rect 2332 1756 2340 1764
rect 2364 1756 2372 1764
rect 2524 1756 2532 1764
rect 2636 1756 2644 1764
rect 460 1736 468 1744
rect 476 1736 484 1744
rect 588 1736 596 1744
rect 12 1716 20 1724
rect 108 1716 116 1724
rect 172 1716 180 1724
rect 316 1716 324 1724
rect 364 1716 372 1724
rect 524 1716 532 1724
rect 588 1716 596 1724
rect 620 1736 628 1744
rect 684 1736 692 1744
rect 716 1736 724 1744
rect 812 1736 820 1744
rect 1052 1736 1060 1744
rect 1372 1736 1380 1744
rect 1484 1736 1492 1744
rect 1676 1736 1684 1744
rect 1692 1736 1700 1744
rect 1740 1736 1748 1744
rect 1900 1736 1908 1744
rect 1948 1736 1956 1744
rect 2252 1736 2260 1744
rect 2380 1736 2388 1744
rect 668 1716 676 1724
rect 732 1716 740 1724
rect 748 1716 756 1724
rect 764 1716 772 1724
rect 876 1716 884 1724
rect 1020 1716 1028 1724
rect 1036 1716 1044 1724
rect 1180 1716 1188 1724
rect 1244 1716 1252 1724
rect 1324 1716 1332 1724
rect 2428 1736 2436 1744
rect 2460 1736 2468 1744
rect 188 1696 196 1704
rect 204 1696 212 1704
rect 492 1696 500 1704
rect 684 1696 692 1704
rect 1596 1716 1604 1724
rect 1660 1716 1668 1724
rect 1804 1716 1812 1724
rect 1900 1716 1908 1724
rect 1996 1716 2004 1724
rect 2044 1716 2052 1724
rect 2220 1716 2228 1724
rect 2284 1716 2292 1724
rect 2412 1716 2420 1724
rect 2428 1716 2436 1724
rect 2476 1716 2484 1724
rect 2556 1716 2564 1724
rect 2604 1716 2612 1724
rect 2876 1756 2884 1764
rect 3372 1756 3380 1764
rect 3404 1756 3412 1764
rect 3420 1756 3428 1764
rect 3500 1756 3508 1764
rect 3740 1756 3748 1764
rect 3804 1756 3812 1764
rect 4380 1756 4388 1764
rect 4764 1756 4772 1764
rect 4924 1756 4932 1764
rect 4988 1756 4996 1764
rect 5068 1756 5076 1764
rect 5724 1756 5732 1764
rect 6012 1756 6020 1764
rect 2860 1736 2868 1744
rect 2924 1736 2932 1744
rect 2940 1736 2948 1744
rect 3308 1736 3316 1744
rect 3436 1736 3444 1744
rect 3500 1736 3508 1744
rect 3532 1736 3540 1744
rect 3564 1736 3572 1744
rect 3628 1736 3636 1744
rect 3692 1736 3700 1744
rect 2668 1716 2676 1724
rect 2700 1716 2708 1724
rect 2828 1716 2836 1724
rect 3228 1716 3236 1724
rect 3292 1716 3300 1724
rect 3564 1716 3572 1724
rect 3580 1716 3588 1724
rect 3644 1716 3652 1724
rect 3692 1716 3700 1724
rect 3900 1736 3908 1744
rect 4108 1736 4116 1744
rect 4204 1736 4212 1744
rect 4332 1736 4340 1744
rect 4700 1736 4708 1744
rect 4860 1736 4868 1744
rect 4908 1736 4916 1744
rect 4956 1736 4964 1744
rect 5020 1736 5028 1744
rect 5132 1736 5140 1744
rect 5148 1736 5156 1744
rect 5260 1736 5268 1744
rect 5436 1736 5444 1744
rect 5468 1736 5476 1744
rect 5548 1736 5556 1744
rect 5580 1736 5588 1744
rect 5628 1736 5636 1744
rect 5644 1736 5652 1744
rect 5708 1736 5716 1744
rect 5788 1736 5796 1744
rect 5820 1736 5828 1744
rect 3836 1716 3844 1724
rect 3884 1716 3892 1724
rect 3964 1718 3972 1726
rect 4188 1716 4196 1724
rect 4268 1716 4276 1724
rect 4284 1716 4292 1724
rect 4524 1716 4532 1724
rect 4716 1716 4724 1724
rect 156 1676 164 1684
rect 1468 1676 1476 1684
rect 1516 1676 1524 1684
rect 1932 1696 1940 1704
rect 1980 1696 1988 1704
rect 2156 1696 2164 1704
rect 2220 1696 2228 1704
rect 2316 1696 2324 1704
rect 2412 1696 2420 1704
rect 2620 1696 2628 1704
rect 2732 1696 2740 1704
rect 2844 1696 2852 1704
rect 2892 1696 2900 1704
rect 2972 1696 2980 1704
rect 3612 1696 3620 1704
rect 3724 1696 3732 1704
rect 3852 1696 3860 1704
rect 4232 1696 4240 1704
rect 4252 1696 4260 1704
rect 4444 1696 4452 1704
rect 4716 1696 4724 1704
rect 4796 1716 4804 1724
rect 4860 1716 4868 1724
rect 4972 1716 4980 1724
rect 5036 1716 5044 1724
rect 5068 1716 5076 1724
rect 5132 1716 5140 1724
rect 4812 1696 4820 1704
rect 4876 1696 4884 1704
rect 5196 1696 5204 1704
rect 5260 1716 5268 1724
rect 5388 1716 5396 1724
rect 5484 1716 5492 1724
rect 5244 1696 5252 1704
rect 5516 1696 5524 1704
rect 5580 1716 5588 1724
rect 5660 1716 5668 1724
rect 5692 1716 5700 1724
rect 5756 1716 5764 1724
rect 5836 1716 5844 1724
rect 6012 1718 6020 1726
rect 6140 1716 6148 1724
rect 6188 1716 6196 1724
rect 5596 1696 5604 1704
rect 5804 1696 5812 1704
rect 5868 1696 5876 1704
rect 1820 1676 1828 1684
rect 2428 1676 2436 1684
rect 2556 1676 2564 1684
rect 2588 1676 2596 1684
rect 2812 1676 2820 1684
rect 3276 1676 3284 1684
rect 4124 1676 4132 1684
rect 5276 1676 5284 1684
rect 172 1656 180 1664
rect 2748 1656 2756 1664
rect 2908 1656 2916 1664
rect 3884 1656 3892 1664
rect 4652 1656 4660 1664
rect 5836 1656 5844 1664
rect 1260 1636 1268 1644
rect 1564 1636 1572 1644
rect 1596 1636 1604 1644
rect 1804 1636 1812 1644
rect 2284 1636 2292 1644
rect 2604 1636 2612 1644
rect 2700 1636 2708 1644
rect 3580 1636 3588 1644
rect 3756 1636 3764 1644
rect 4412 1636 4420 1644
rect 4844 1636 4852 1644
rect 5884 1636 5892 1644
rect 1577 1606 1585 1614
rect 1587 1606 1595 1614
rect 1597 1606 1605 1614
rect 1607 1606 1615 1614
rect 4665 1606 4673 1614
rect 4675 1606 4683 1614
rect 4685 1606 4693 1614
rect 4695 1606 4703 1614
rect 364 1576 372 1584
rect 428 1576 436 1584
rect 668 1576 676 1584
rect 1308 1576 1316 1584
rect 1388 1576 1396 1584
rect 1692 1576 1700 1584
rect 1756 1576 1764 1584
rect 1996 1576 2004 1584
rect 2236 1576 2244 1584
rect 2268 1576 2276 1584
rect 2380 1576 2388 1584
rect 2860 1576 2868 1584
rect 3180 1576 3188 1584
rect 4044 1576 4052 1584
rect 4876 1576 4884 1584
rect 4908 1576 4916 1584
rect 5084 1576 5092 1584
rect 5452 1576 5460 1584
rect 5468 1576 5476 1584
rect 5804 1576 5812 1584
rect 316 1556 324 1564
rect 92 1536 100 1544
rect 620 1536 628 1544
rect 1020 1536 1028 1544
rect 1132 1536 1140 1544
rect 1196 1536 1204 1544
rect 1276 1536 1284 1544
rect 1980 1536 1988 1544
rect 2476 1536 2484 1544
rect 2556 1556 2564 1564
rect 6108 1556 6116 1564
rect 2508 1536 2516 1544
rect 2588 1536 2596 1544
rect 2988 1536 2996 1544
rect 3500 1536 3508 1544
rect 3724 1536 3732 1544
rect 4252 1536 4260 1544
rect 4380 1536 4388 1544
rect 4636 1536 4644 1544
rect 4668 1536 4676 1544
rect 4732 1536 4740 1544
rect 5964 1536 5972 1544
rect 6012 1536 6020 1544
rect 12 1516 20 1524
rect 44 1516 52 1524
rect 220 1496 228 1504
rect 396 1496 404 1504
rect 428 1496 436 1504
rect 540 1516 548 1524
rect 844 1516 852 1524
rect 876 1516 884 1524
rect 940 1516 948 1524
rect 988 1516 996 1524
rect 1052 1516 1060 1524
rect 1164 1516 1172 1524
rect 1228 1516 1236 1524
rect 1244 1516 1252 1524
rect 1420 1516 1428 1524
rect 1612 1516 1620 1524
rect 60 1476 68 1484
rect 268 1476 276 1484
rect 300 1476 308 1484
rect 332 1476 340 1484
rect 412 1476 420 1484
rect 524 1496 532 1504
rect 604 1496 612 1504
rect 684 1496 692 1504
rect 700 1496 708 1504
rect 572 1476 580 1484
rect 92 1456 100 1464
rect 652 1456 660 1464
rect 732 1496 740 1504
rect 748 1496 756 1504
rect 796 1496 804 1504
rect 844 1496 852 1504
rect 1036 1496 1044 1504
rect 1084 1496 1092 1504
rect 1212 1496 1220 1504
rect 1260 1496 1268 1504
rect 1340 1496 1348 1504
rect 1388 1496 1396 1504
rect 732 1476 740 1484
rect 892 1476 900 1484
rect 956 1476 964 1484
rect 1068 1476 1076 1484
rect 1132 1476 1140 1484
rect 1148 1476 1156 1484
rect 1372 1476 1380 1484
rect 1436 1476 1444 1484
rect 1484 1496 1492 1504
rect 1484 1476 1492 1484
rect 1548 1476 1556 1484
rect 1676 1496 1684 1504
rect 1772 1516 1780 1524
rect 2012 1516 2020 1524
rect 2300 1516 2308 1524
rect 2444 1516 2452 1524
rect 2508 1516 2516 1524
rect 2604 1516 2612 1524
rect 2764 1516 2772 1524
rect 2924 1516 2932 1524
rect 2972 1516 2980 1524
rect 3020 1516 3028 1524
rect 3228 1516 3236 1524
rect 3948 1516 3956 1524
rect 1804 1496 1812 1504
rect 1836 1496 1844 1504
rect 1996 1496 2004 1504
rect 2156 1496 2164 1504
rect 2188 1496 2196 1504
rect 2252 1496 2260 1504
rect 2268 1496 2276 1504
rect 2332 1496 2340 1504
rect 2396 1496 2404 1504
rect 2412 1496 2420 1504
rect 2492 1496 2500 1504
rect 2556 1496 2564 1504
rect 2588 1496 2596 1504
rect 2636 1496 2644 1504
rect 2668 1496 2676 1504
rect 2684 1496 2692 1504
rect 2796 1496 2804 1504
rect 2876 1496 2884 1504
rect 2892 1496 2900 1504
rect 2940 1496 2948 1504
rect 3004 1496 3012 1504
rect 3116 1496 3124 1504
rect 3148 1496 3156 1504
rect 3260 1496 3268 1504
rect 3340 1494 3348 1502
rect 3612 1496 3620 1504
rect 3692 1496 3700 1504
rect 3708 1496 3716 1504
rect 4124 1516 4132 1524
rect 4156 1516 4164 1524
rect 4684 1516 4692 1524
rect 4764 1516 4772 1524
rect 3852 1494 3860 1502
rect 4060 1496 4068 1504
rect 4156 1496 4164 1504
rect 4252 1496 4260 1504
rect 4284 1496 4292 1504
rect 4508 1496 4516 1504
rect 4956 1516 4964 1524
rect 5276 1516 5284 1524
rect 5308 1516 5316 1524
rect 5340 1516 5348 1524
rect 5772 1516 5780 1524
rect 5836 1516 5844 1524
rect 5944 1516 5952 1524
rect 5980 1516 5988 1524
rect 6044 1516 6052 1524
rect 4812 1496 4820 1504
rect 4876 1496 4884 1504
rect 4940 1496 4948 1504
rect 5020 1496 5028 1504
rect 5212 1494 5220 1502
rect 5308 1496 5316 1504
rect 5324 1496 5332 1504
rect 5532 1496 5540 1504
rect 5548 1496 5556 1504
rect 5660 1496 5668 1504
rect 1676 1476 1684 1484
rect 1740 1476 1748 1484
rect 2140 1476 2148 1484
rect 2316 1476 2324 1484
rect 2348 1476 2356 1484
rect 2396 1476 2404 1484
rect 2428 1476 2436 1484
rect 2636 1476 2644 1484
rect 2812 1476 2820 1484
rect 2860 1476 2868 1484
rect 3276 1476 3284 1484
rect 3628 1476 3636 1484
rect 3644 1476 3652 1484
rect 3916 1476 3924 1484
rect 3948 1476 3956 1484
rect 4012 1476 4020 1484
rect 4028 1476 4036 1484
rect 4172 1476 4180 1484
rect 4268 1476 4276 1484
rect 4284 1476 4292 1484
rect 4348 1476 4356 1484
rect 4588 1476 4596 1484
rect 4636 1476 4644 1484
rect 4732 1476 4740 1484
rect 4828 1476 4836 1484
rect 4988 1476 4996 1484
rect 5244 1476 5252 1484
rect 5324 1476 5332 1484
rect 5420 1476 5428 1484
rect 5484 1476 5492 1484
rect 5724 1496 5732 1504
rect 5740 1496 5748 1504
rect 5804 1496 5812 1504
rect 5836 1496 5844 1504
rect 5932 1496 5940 1504
rect 6012 1496 6020 1504
rect 6028 1496 6036 1504
rect 6076 1496 6084 1504
rect 6220 1496 6228 1504
rect 5724 1476 5732 1484
rect 5756 1476 5764 1484
rect 5788 1476 5796 1484
rect 5852 1476 5860 1484
rect 5916 1476 5924 1484
rect 6028 1476 6036 1484
rect 6092 1476 6100 1484
rect 6204 1476 6212 1484
rect 828 1456 836 1464
rect 1516 1456 1524 1464
rect 1564 1456 1572 1464
rect 1740 1456 1748 1464
rect 1772 1456 1780 1464
rect 1868 1456 1876 1464
rect 1948 1456 1956 1464
rect 2124 1456 2132 1464
rect 2220 1456 2228 1464
rect 2284 1456 2292 1464
rect 2524 1456 2532 1464
rect 2828 1456 2836 1464
rect 2940 1456 2948 1464
rect 3036 1456 3044 1464
rect 3228 1456 3236 1464
rect 4188 1456 4196 1464
rect 4524 1456 4532 1464
rect 4844 1456 4852 1464
rect 5004 1456 5012 1464
rect 5404 1456 5412 1464
rect 492 1436 500 1444
rect 620 1436 628 1444
rect 780 1436 788 1444
rect 988 1436 996 1444
rect 1292 1436 1300 1444
rect 1564 1436 1572 1444
rect 1900 1436 1908 1444
rect 2588 1436 2596 1444
rect 2668 1436 2676 1444
rect 3084 1436 3092 1444
rect 3100 1436 3108 1444
rect 3468 1436 3476 1444
rect 3564 1436 3572 1444
rect 4044 1436 4052 1444
rect 4092 1436 4100 1444
rect 4396 1436 4404 1444
rect 4780 1436 4788 1444
rect 4908 1436 4916 1444
rect 5052 1436 5060 1444
rect 5900 1436 5908 1444
rect 3113 1406 3121 1414
rect 3123 1406 3131 1414
rect 3133 1406 3141 1414
rect 3143 1406 3151 1414
rect 12 1376 20 1384
rect 204 1376 212 1384
rect 316 1376 324 1384
rect 572 1376 580 1384
rect 636 1376 644 1384
rect 1132 1376 1140 1384
rect 1260 1376 1268 1384
rect 1356 1376 1364 1384
rect 1724 1376 1732 1384
rect 1964 1376 1972 1384
rect 2300 1376 2308 1384
rect 2764 1376 2772 1384
rect 2972 1376 2980 1384
rect 3244 1376 3252 1384
rect 3324 1376 3332 1384
rect 3916 1376 3924 1384
rect 4108 1376 4116 1384
rect 4620 1376 4628 1384
rect 4924 1376 4932 1384
rect 5052 1376 5060 1384
rect 5180 1376 5188 1384
rect 5500 1376 5508 1384
rect 5612 1376 5620 1384
rect 5804 1376 5812 1384
rect 6076 1376 6084 1384
rect 156 1356 164 1364
rect 188 1356 196 1364
rect 332 1356 340 1364
rect 396 1356 404 1364
rect 412 1356 420 1364
rect 444 1356 452 1364
rect 476 1356 484 1364
rect 716 1356 724 1364
rect 1020 1356 1028 1364
rect 1372 1356 1380 1364
rect 1404 1356 1412 1364
rect 1452 1356 1460 1364
rect 1612 1356 1620 1364
rect 1852 1356 1860 1364
rect 1900 1356 1908 1364
rect 2140 1356 2148 1364
rect 2236 1356 2244 1364
rect 2316 1356 2324 1364
rect 2636 1356 2644 1364
rect 3052 1356 3060 1364
rect 3084 1356 3092 1364
rect 3628 1356 3636 1364
rect 3932 1356 3940 1364
rect 5004 1356 5012 1364
rect 5132 1356 5140 1364
rect 5164 1356 5172 1364
rect 6204 1356 6212 1364
rect 44 1336 52 1344
rect 60 1336 68 1344
rect 188 1336 196 1344
rect 316 1336 324 1344
rect 412 1336 420 1344
rect 524 1336 532 1344
rect 588 1336 596 1344
rect 652 1336 660 1344
rect 684 1336 692 1344
rect 748 1336 756 1344
rect 812 1336 820 1344
rect 940 1336 948 1344
rect 972 1336 980 1344
rect 1036 1336 1044 1344
rect 1068 1336 1076 1344
rect 1100 1336 1108 1344
rect 1148 1336 1156 1344
rect 1164 1336 1172 1344
rect 1388 1336 1396 1344
rect 1436 1336 1444 1344
rect 1532 1336 1540 1344
rect 1644 1336 1652 1344
rect 1868 1336 1876 1344
rect 2108 1336 2116 1344
rect 2156 1336 2164 1344
rect 2300 1336 2308 1344
rect 2396 1336 2404 1344
rect 124 1316 132 1324
rect 220 1316 228 1324
rect 300 1316 308 1324
rect 316 1316 324 1324
rect 412 1316 420 1324
rect 652 1316 660 1324
rect 12 1296 20 1304
rect 572 1296 580 1304
rect 956 1316 964 1324
rect 988 1316 996 1324
rect 1084 1316 1092 1324
rect 812 1296 820 1304
rect 1212 1316 1220 1324
rect 1324 1316 1332 1324
rect 1548 1316 1556 1324
rect 1756 1316 1764 1324
rect 1788 1316 1796 1324
rect 2172 1316 2180 1324
rect 2396 1316 2404 1324
rect 2524 1336 2532 1344
rect 2556 1336 2564 1344
rect 2588 1336 2596 1344
rect 2716 1336 2724 1344
rect 2780 1336 2788 1344
rect 2796 1336 2804 1344
rect 2860 1336 2868 1344
rect 2924 1336 2932 1344
rect 2988 1336 2996 1344
rect 3244 1336 3252 1344
rect 3276 1336 3284 1344
rect 3292 1336 3300 1344
rect 3388 1336 3396 1344
rect 3788 1336 3796 1344
rect 4092 1336 4100 1344
rect 4300 1336 4308 1344
rect 4348 1336 4356 1344
rect 4412 1336 4420 1344
rect 4732 1336 4740 1344
rect 4828 1336 4836 1344
rect 4908 1336 4916 1344
rect 4972 1336 4980 1344
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 5292 1336 5300 1344
rect 5420 1336 5428 1344
rect 5548 1336 5556 1344
rect 5596 1336 5604 1344
rect 5964 1336 5972 1344
rect 6012 1336 6020 1344
rect 6044 1336 6052 1344
rect 2428 1316 2436 1324
rect 2636 1316 2644 1324
rect 2732 1316 2740 1324
rect 2764 1316 2772 1324
rect 2796 1316 2804 1324
rect 2812 1316 2820 1324
rect 2876 1316 2884 1324
rect 3004 1316 3012 1324
rect 3180 1316 3188 1324
rect 3532 1318 3540 1326
rect 3596 1316 3604 1324
rect 3676 1316 3684 1324
rect 3804 1316 3812 1324
rect 3964 1316 3972 1324
rect 4028 1316 4036 1324
rect 4060 1316 4068 1324
rect 4076 1316 4084 1324
rect 4172 1316 4180 1324
rect 4220 1316 4228 1324
rect 4348 1316 4356 1324
rect 4396 1316 4404 1324
rect 4476 1318 4484 1326
rect 4524 1316 4532 1324
rect 4764 1316 4772 1324
rect 4892 1316 4900 1324
rect 4956 1316 4964 1324
rect 5084 1316 5092 1324
rect 5100 1316 5108 1324
rect 5132 1316 5140 1324
rect 5276 1316 5284 1324
rect 5372 1316 5380 1324
rect 5452 1316 5460 1324
rect 1212 1296 1220 1304
rect 1468 1296 1476 1304
rect 1484 1296 1492 1304
rect 1516 1296 1524 1304
rect 1724 1296 1732 1304
rect 2460 1296 2468 1304
rect 2652 1296 2660 1304
rect 2972 1296 2980 1304
rect 3692 1296 3700 1304
rect 3724 1296 3732 1304
rect 3980 1296 3988 1304
rect 4012 1296 4020 1304
rect 4316 1296 4324 1304
rect 4332 1296 4340 1304
rect 4396 1296 4404 1304
rect 4892 1296 4900 1304
rect 4924 1296 4932 1304
rect 5020 1296 5028 1304
rect 5484 1296 5492 1304
rect 5532 1316 5540 1324
rect 5676 1316 5684 1324
rect 5724 1316 5732 1324
rect 5916 1316 5924 1324
rect 5996 1316 6004 1324
rect 6028 1316 6036 1324
rect 6060 1316 6068 1324
rect 6188 1316 6196 1324
rect 5564 1296 5572 1304
rect 1324 1276 1332 1284
rect 2684 1276 2692 1284
rect 3036 1276 3044 1284
rect 6108 1276 6116 1284
rect 5580 1256 5588 1264
rect 732 1236 740 1244
rect 828 1236 836 1244
rect 1756 1236 1764 1244
rect 2012 1236 2020 1244
rect 2124 1236 2132 1244
rect 2428 1236 2436 1244
rect 2604 1236 2612 1244
rect 2668 1236 2676 1244
rect 3052 1236 3060 1244
rect 3116 1236 3124 1244
rect 3212 1236 3220 1244
rect 3596 1236 3604 1244
rect 5100 1236 5108 1244
rect 1577 1206 1585 1214
rect 1587 1206 1595 1214
rect 1597 1206 1605 1214
rect 1607 1206 1615 1214
rect 4665 1206 4673 1214
rect 4675 1206 4683 1214
rect 4685 1206 4693 1214
rect 4695 1206 4703 1214
rect 44 1176 52 1184
rect 156 1176 164 1184
rect 300 1176 308 1184
rect 572 1176 580 1184
rect 924 1176 932 1184
rect 1068 1176 1076 1184
rect 1276 1176 1284 1184
rect 1356 1176 1364 1184
rect 1836 1176 1844 1184
rect 1868 1176 1876 1184
rect 2076 1176 2084 1184
rect 2380 1176 2388 1184
rect 2652 1176 2660 1184
rect 3180 1176 3188 1184
rect 3580 1176 3588 1184
rect 3916 1176 3924 1184
rect 4140 1176 4148 1184
rect 4252 1176 4260 1184
rect 4908 1176 4916 1184
rect 4972 1176 4980 1184
rect 5020 1176 5028 1184
rect 5148 1176 5156 1184
rect 5180 1176 5188 1184
rect 5308 1176 5316 1184
rect 5516 1176 5524 1184
rect 5580 1176 5588 1184
rect 5676 1176 5684 1184
rect 5724 1176 5732 1184
rect 5868 1176 5876 1184
rect 6012 1176 6020 1184
rect 6140 1176 6148 1184
rect 6220 1176 6228 1184
rect 1692 1156 1700 1164
rect 2716 1156 2724 1164
rect 3612 1156 3620 1164
rect 4284 1156 4292 1164
rect 508 1136 516 1144
rect 556 1136 564 1144
rect 668 1136 676 1144
rect 684 1136 692 1144
rect 732 1136 740 1144
rect 812 1136 820 1144
rect 988 1136 996 1144
rect 1132 1136 1140 1144
rect 1292 1136 1300 1144
rect 4124 1136 4132 1144
rect 4316 1136 4324 1144
rect 5132 1136 5140 1144
rect 524 1116 532 1124
rect 588 1116 596 1124
rect 636 1116 644 1124
rect 700 1116 708 1124
rect 764 1116 772 1124
rect 12 1096 20 1104
rect 124 1096 132 1104
rect 172 1096 180 1104
rect 204 1096 212 1104
rect 220 1096 228 1104
rect 316 1096 324 1104
rect 460 1096 468 1104
rect 492 1096 500 1104
rect 572 1096 580 1104
rect 684 1096 692 1104
rect 748 1096 756 1104
rect 780 1096 788 1104
rect 828 1096 836 1104
rect 908 1116 916 1124
rect 940 1116 948 1124
rect 988 1116 996 1124
rect 1036 1116 1044 1124
rect 908 1096 916 1104
rect 1196 1116 1204 1124
rect 1260 1116 1268 1124
rect 1340 1116 1348 1124
rect 1484 1116 1492 1124
rect 1532 1116 1540 1124
rect 1548 1116 1556 1124
rect 2124 1116 2132 1124
rect 2396 1116 2404 1124
rect 2444 1116 2452 1124
rect 3116 1116 3124 1124
rect 3404 1116 3412 1124
rect 428 1076 436 1084
rect 604 1076 612 1084
rect 844 1076 852 1084
rect 940 1076 948 1084
rect 988 1076 996 1084
rect 1036 1076 1044 1084
rect 1084 1076 1092 1084
rect 1132 1076 1140 1084
rect 1164 1096 1172 1104
rect 1244 1096 1252 1104
rect 1308 1096 1316 1104
rect 1436 1096 1444 1104
rect 1484 1096 1492 1104
rect 1708 1096 1716 1104
rect 1884 1096 1892 1104
rect 1900 1096 1908 1104
rect 1980 1096 1988 1104
rect 2172 1096 2180 1104
rect 2220 1096 2228 1104
rect 2284 1096 2292 1104
rect 2412 1096 2420 1104
rect 2476 1096 2484 1104
rect 2524 1096 2532 1104
rect 2556 1096 2564 1104
rect 2796 1096 2804 1104
rect 2876 1096 2884 1104
rect 2924 1096 2932 1104
rect 2972 1096 2980 1104
rect 3020 1096 3028 1104
rect 3084 1096 3092 1104
rect 3116 1096 3124 1104
rect 3164 1096 3172 1104
rect 3292 1096 3300 1104
rect 4732 1116 4740 1124
rect 4796 1116 4804 1124
rect 4940 1116 4948 1124
rect 5052 1116 5060 1124
rect 5340 1116 5348 1124
rect 3452 1096 3460 1104
rect 3500 1096 3508 1104
rect 3756 1094 3764 1102
rect 3820 1096 3828 1104
rect 3852 1096 3860 1104
rect 3868 1096 3876 1104
rect 3996 1096 4004 1104
rect 4044 1096 4052 1104
rect 4220 1096 4228 1104
rect 4348 1096 4356 1104
rect 4364 1096 4372 1104
rect 1340 1076 1348 1084
rect 1516 1076 1524 1084
rect 1548 1076 1556 1084
rect 1996 1076 2004 1084
rect 2012 1076 2020 1084
rect 2156 1076 2164 1084
rect 2252 1076 2260 1084
rect 2364 1076 2372 1084
rect 2444 1076 2452 1084
rect 2508 1076 2516 1084
rect 2620 1076 2628 1084
rect 2764 1076 2772 1084
rect 2828 1076 2836 1084
rect 2844 1076 2852 1084
rect 3068 1076 3076 1084
rect 3308 1076 3316 1084
rect 3372 1076 3380 1084
rect 3420 1076 3428 1084
rect 3468 1076 3476 1084
rect 3724 1076 3732 1084
rect 3820 1076 3828 1084
rect 3884 1076 3892 1084
rect 4172 1076 4180 1084
rect 76 1056 84 1064
rect 124 1056 132 1064
rect 172 1056 180 1064
rect 268 1056 276 1064
rect 316 1056 324 1064
rect 380 1056 388 1064
rect 428 1056 436 1064
rect 1708 1056 1716 1064
rect 1740 1056 1748 1064
rect 1804 1056 1812 1064
rect 1852 1056 1860 1064
rect 2204 1056 2212 1064
rect 2252 1056 2260 1064
rect 2556 1056 2564 1064
rect 2636 1056 2644 1064
rect 2828 1056 2836 1064
rect 2860 1056 2868 1064
rect 3052 1056 3060 1064
rect 3516 1056 3524 1064
rect 3548 1056 3556 1064
rect 3564 1056 3572 1064
rect 3596 1056 3604 1064
rect 3900 1056 3908 1064
rect 4124 1056 4132 1064
rect 4204 1056 4212 1064
rect 4300 1056 4308 1064
rect 4476 1096 4484 1104
rect 4524 1096 4532 1104
rect 4620 1096 4628 1104
rect 4652 1096 4660 1104
rect 4828 1096 4836 1104
rect 4844 1096 4852 1104
rect 4924 1096 4932 1104
rect 4988 1096 4996 1104
rect 5100 1096 5108 1104
rect 5148 1096 5156 1104
rect 5212 1096 5220 1104
rect 5292 1096 5300 1104
rect 5372 1096 5380 1104
rect 5644 1116 5652 1124
rect 5756 1116 5764 1124
rect 5820 1116 5828 1124
rect 5836 1116 5844 1124
rect 6252 1116 6260 1124
rect 5436 1096 5444 1104
rect 5468 1096 5476 1104
rect 5532 1096 5540 1104
rect 5596 1096 5604 1104
rect 5708 1096 5716 1104
rect 5724 1096 5732 1104
rect 5788 1096 5796 1104
rect 5804 1096 5812 1104
rect 5884 1096 5892 1104
rect 5900 1096 5908 1104
rect 6028 1096 6036 1104
rect 6092 1096 6100 1104
rect 6220 1096 6228 1104
rect 4684 1076 4692 1084
rect 4780 1076 4788 1084
rect 4844 1076 4852 1084
rect 4876 1076 4884 1084
rect 4924 1076 4932 1084
rect 4988 1076 4996 1084
rect 5100 1076 5108 1084
rect 5324 1076 5332 1084
rect 5372 1076 5380 1084
rect 5388 1076 5396 1084
rect 5548 1076 5556 1084
rect 5596 1076 5604 1084
rect 5612 1076 5620 1084
rect 5708 1076 5716 1084
rect 5772 1076 5780 1084
rect 5884 1076 5892 1084
rect 6044 1076 6052 1084
rect 6076 1076 6084 1084
rect 6172 1076 6180 1084
rect 6188 1076 6196 1084
rect 4380 1056 4388 1064
rect 4396 1056 4404 1064
rect 5004 1056 5012 1064
rect 5244 1056 5252 1064
rect 5324 1056 5332 1064
rect 5436 1056 5444 1064
rect 5484 1056 5492 1064
rect 5628 1056 5636 1064
rect 5932 1056 5940 1064
rect 5996 1056 6004 1064
rect 6124 1056 6132 1064
rect 6188 1056 6196 1064
rect 92 1036 100 1044
rect 332 1036 340 1044
rect 636 1036 644 1044
rect 1020 1036 1028 1044
rect 1100 1036 1108 1044
rect 1228 1036 1236 1044
rect 1788 1036 1796 1044
rect 1916 1036 1924 1044
rect 2060 1036 2068 1044
rect 2316 1036 2324 1044
rect 2732 1036 2740 1044
rect 3004 1036 3012 1044
rect 3164 1036 3172 1044
rect 3484 1036 3492 1044
rect 3628 1036 3636 1044
rect 4188 1036 4196 1044
rect 4588 1036 4596 1044
rect 4652 1036 4660 1044
rect 4700 1036 4708 1044
rect 5180 1036 5188 1044
rect 5276 1036 5284 1044
rect 5500 1036 5508 1044
rect 6044 1036 6052 1044
rect 3113 1006 3121 1014
rect 3123 1006 3131 1014
rect 3133 1006 3141 1014
rect 3143 1006 3151 1014
rect 44 976 52 984
rect 76 976 84 984
rect 172 976 180 984
rect 204 976 212 984
rect 348 976 356 984
rect 444 976 452 984
rect 796 976 804 984
rect 908 976 916 984
rect 1084 976 1092 984
rect 1180 976 1188 984
rect 2076 976 2084 984
rect 2748 976 2756 984
rect 3020 976 3028 984
rect 3500 976 3508 984
rect 3612 976 3620 984
rect 3884 976 3892 984
rect 3916 976 3924 984
rect 4124 976 4132 984
rect 4364 976 4372 984
rect 4476 976 4484 984
rect 4780 976 4788 984
rect 5132 976 5140 984
rect 5356 976 5364 984
rect 5532 976 5540 984
rect 5564 976 5572 984
rect 5756 976 5764 984
rect 5948 976 5956 984
rect 6028 976 6036 984
rect 6044 976 6052 984
rect 140 956 148 964
rect 268 956 276 964
rect 364 956 372 964
rect 396 956 404 964
rect 492 956 500 964
rect 524 956 532 964
rect 12 936 20 944
rect 60 936 68 944
rect 92 936 100 944
rect 188 936 196 944
rect 252 936 260 944
rect 300 936 308 944
rect 476 936 484 944
rect 924 956 932 964
rect 956 956 964 964
rect 1004 956 1012 964
rect 1020 956 1028 964
rect 1228 956 1236 964
rect 1580 956 1588 964
rect 1596 956 1604 964
rect 1644 956 1652 964
rect 1980 956 1988 964
rect 700 936 708 944
rect 764 936 772 944
rect 860 936 868 944
rect 876 936 884 944
rect 908 936 916 944
rect 316 916 324 924
rect 412 916 420 924
rect 492 916 500 924
rect 652 916 660 924
rect 700 916 708 924
rect 828 916 836 924
rect 988 936 996 944
rect 1020 936 1028 944
rect 1052 936 1060 944
rect 1116 936 1124 944
rect 1164 936 1172 944
rect 1196 936 1204 944
rect 1340 936 1348 944
rect 1452 936 1460 944
rect 1532 936 1540 944
rect 1740 936 1748 944
rect 1772 936 1780 944
rect 1836 936 1844 944
rect 2060 956 2068 964
rect 2108 956 2116 964
rect 2348 956 2356 964
rect 2380 956 2388 964
rect 2460 956 2468 964
rect 2556 956 2564 964
rect 2588 956 2596 964
rect 2604 956 2612 964
rect 2844 956 2852 964
rect 2860 956 2868 964
rect 3276 956 3284 964
rect 3372 956 3380 964
rect 3596 956 3604 964
rect 3900 956 3908 964
rect 4044 956 4052 964
rect 4348 956 4356 964
rect 4892 956 4900 964
rect 4924 956 4932 964
rect 5116 956 5124 964
rect 5212 956 5220 964
rect 5436 956 5444 964
rect 5628 956 5636 964
rect 5692 956 5700 964
rect 5740 956 5748 964
rect 5836 956 5844 964
rect 5900 956 5908 964
rect 5932 956 5940 964
rect 5964 956 5972 964
rect 2060 936 2068 944
rect 2140 936 2148 944
rect 2220 936 2228 944
rect 2332 936 2340 944
rect 2460 936 2468 944
rect 2492 936 2500 944
rect 2588 936 2596 944
rect 2876 936 2884 944
rect 2956 936 2964 944
rect 2988 936 2996 944
rect 3292 936 3300 944
rect 3516 936 3524 944
rect 3564 936 3572 944
rect 3724 936 3732 944
rect 3804 936 3812 944
rect 3836 936 3844 944
rect 4252 936 4260 944
rect 4412 936 4420 944
rect 4604 936 4612 944
rect 4716 936 4724 944
rect 4748 936 4756 944
rect 4828 936 4836 944
rect 4988 936 4996 944
rect 5100 936 5108 944
rect 5228 936 5236 944
rect 972 916 980 924
rect 1276 916 1284 924
rect 1612 916 1620 924
rect 1660 916 1668 924
rect 1756 916 1764 924
rect 1836 916 1844 924
rect 1932 916 1940 924
rect 2092 916 2100 924
rect 2172 916 2180 924
rect 2220 916 2228 924
rect 2236 916 2244 924
rect 2268 916 2276 924
rect 2348 916 2356 924
rect 2492 916 2500 924
rect 2540 916 2548 924
rect 2700 916 2708 924
rect 2732 916 2740 924
rect 2844 916 2852 924
rect 2892 916 2900 924
rect 60 896 68 904
rect 92 896 100 904
rect 156 896 164 904
rect 204 896 212 904
rect 236 896 244 904
rect 540 896 548 904
rect 620 896 628 904
rect 748 896 756 904
rect 796 896 804 904
rect 812 896 820 904
rect 908 896 916 904
rect 1164 896 1172 904
rect 1292 896 1300 904
rect 1484 896 1492 904
rect 1516 896 1524 904
rect 1708 896 1716 904
rect 1932 896 1940 904
rect 2204 896 2212 904
rect 2284 896 2292 904
rect 2540 896 2548 904
rect 2716 896 2724 904
rect 2924 896 2932 904
rect 2972 916 2980 924
rect 3020 916 3028 924
rect 3084 916 3092 924
rect 3212 916 3220 924
rect 3244 916 3252 924
rect 3308 916 3316 924
rect 3388 916 3396 924
rect 3564 916 3572 924
rect 3740 918 3748 926
rect 3820 916 3828 924
rect 4044 918 4052 926
rect 4156 916 4164 924
rect 4236 916 4244 924
rect 4268 916 4276 924
rect 4316 916 4324 924
rect 4572 916 4580 924
rect 4732 916 4740 924
rect 4972 916 4980 924
rect 5020 916 5028 924
rect 5052 916 5060 924
rect 5148 916 5156 924
rect 5180 916 5188 924
rect 5228 916 5236 924
rect 5276 916 5284 924
rect 5404 936 5412 944
rect 5436 936 5444 944
rect 5500 936 5508 944
rect 5516 936 5524 944
rect 5964 936 5972 944
rect 5980 936 5988 944
rect 6140 936 6148 944
rect 6236 936 6244 944
rect 5356 916 5364 924
rect 5468 916 5476 924
rect 3068 896 3076 904
rect 3228 896 3236 904
rect 3516 896 3524 904
rect 3852 896 3860 904
rect 4140 896 4148 904
rect 4364 896 4372 904
rect 4492 896 4500 904
rect 4540 896 4548 904
rect 4780 896 4788 904
rect 4876 896 4884 904
rect 4940 896 4948 904
rect 5068 896 5076 904
rect 5212 896 5220 904
rect 5276 896 5284 904
rect 5292 896 5300 904
rect 5356 896 5364 904
rect 5564 916 5572 924
rect 5596 916 5604 924
rect 5724 916 5732 924
rect 5788 916 5796 924
rect 5804 916 5812 924
rect 5932 916 5940 924
rect 5980 916 5988 924
rect 5996 916 6004 924
rect 6172 918 6180 926
rect 6252 916 6260 924
rect 5564 896 5572 904
rect 5628 896 5636 904
rect 6028 896 6036 904
rect 6284 896 6292 904
rect 44 876 52 884
rect 396 876 404 884
rect 604 876 612 884
rect 620 876 628 884
rect 1212 876 1220 884
rect 1260 876 1268 884
rect 1292 876 1300 884
rect 1340 876 1348 884
rect 1948 876 1956 884
rect 3004 876 3012 884
rect 3100 876 3108 884
rect 3196 876 3204 884
rect 4188 876 4196 884
rect 5244 876 5252 884
rect 5436 876 5444 884
rect 6300 876 6308 884
rect 1372 856 1380 864
rect 2028 856 2036 864
rect 2428 856 2436 864
rect 3084 856 3092 864
rect 5884 856 5892 864
rect 428 836 436 844
rect 716 836 724 844
rect 1436 836 1444 844
rect 1468 836 1476 844
rect 1676 836 1684 844
rect 1820 836 1828 844
rect 1932 836 1940 844
rect 2092 836 2100 844
rect 2236 836 2244 844
rect 2652 836 2660 844
rect 2796 836 2804 844
rect 3212 836 3220 844
rect 4204 836 4212 844
rect 4508 836 4516 844
rect 4572 836 4580 844
rect 1577 806 1585 814
rect 1587 806 1595 814
rect 1597 806 1605 814
rect 1607 806 1615 814
rect 4665 806 4673 814
rect 4675 806 4683 814
rect 4685 806 4693 814
rect 4695 806 4703 814
rect 156 776 164 784
rect 188 776 196 784
rect 236 776 244 784
rect 252 776 260 784
rect 332 776 340 784
rect 508 776 516 784
rect 764 776 772 784
rect 844 776 852 784
rect 2844 776 2852 784
rect 3820 776 3828 784
rect 3996 776 4004 784
rect 4044 776 4052 784
rect 4220 776 4228 784
rect 4588 776 4596 784
rect 4620 776 4628 784
rect 4828 776 4836 784
rect 4860 776 4868 784
rect 5068 776 5076 784
rect 5100 776 5108 784
rect 5148 776 5156 784
rect 5228 776 5236 784
rect 5356 776 5364 784
rect 5468 776 5476 784
rect 5692 776 5700 784
rect 5884 776 5892 784
rect 5964 776 5972 784
rect 6092 776 6100 784
rect 6284 776 6292 784
rect 3612 756 3620 764
rect 60 736 68 744
rect 860 736 868 744
rect 956 736 964 744
rect 540 716 548 724
rect 636 716 644 724
rect 668 716 676 724
rect 684 716 692 724
rect 812 716 820 724
rect 828 716 836 724
rect 44 696 52 704
rect 92 696 100 704
rect 348 696 356 704
rect 492 696 500 704
rect 732 696 740 704
rect 844 696 852 704
rect 1084 736 1092 744
rect 1436 736 1444 744
rect 1484 736 1492 744
rect 1644 736 1652 744
rect 3084 736 3092 744
rect 3484 736 3492 744
rect 4060 736 4068 744
rect 4108 736 4116 744
rect 988 716 996 724
rect 1004 716 1012 724
rect 1116 716 1124 724
rect 1164 716 1172 724
rect 1244 716 1252 724
rect 1052 696 1060 704
rect 1100 696 1108 704
rect 1292 696 1300 704
rect 1372 696 1380 704
rect 1724 716 1732 724
rect 1788 716 1796 724
rect 2028 716 2036 724
rect 1756 696 1764 704
rect 1820 696 1828 704
rect 1932 696 1940 704
rect 2156 716 2164 724
rect 2268 716 2276 724
rect 2312 716 2320 724
rect 2332 716 2340 724
rect 2460 716 2468 724
rect 2076 696 2084 704
rect 2124 696 2132 704
rect 2204 696 2212 704
rect 2268 696 2276 704
rect 2396 696 2404 704
rect 2716 716 2724 724
rect 2780 716 2788 724
rect 2904 716 2912 724
rect 2924 716 2932 724
rect 3036 716 3044 724
rect 3132 716 3140 724
rect 3260 716 3268 724
rect 3308 716 3316 724
rect 3372 716 3380 724
rect 2508 696 2516 704
rect 2524 696 2532 704
rect 2572 696 2580 704
rect 2588 696 2596 704
rect 2668 696 2676 704
rect 2700 696 2708 704
rect 2764 696 2772 704
rect 2860 696 2868 704
rect 2940 696 2948 704
rect 2988 696 2996 704
rect 3100 696 3108 704
rect 3180 696 3188 704
rect 3324 696 3332 704
rect 3388 696 3396 704
rect 3404 696 3412 704
rect 3468 696 3476 704
rect 412 676 420 684
rect 444 676 452 684
rect 572 676 580 684
rect 588 676 596 684
rect 620 676 628 684
rect 716 676 724 684
rect 780 676 788 684
rect 892 676 900 684
rect 956 676 964 684
rect 1052 676 1060 684
rect 1132 676 1140 684
rect 1196 676 1204 684
rect 1244 676 1252 684
rect 1276 676 1284 684
rect 1324 676 1332 684
rect 1372 676 1380 684
rect 1420 676 1428 684
rect 1532 676 1540 684
rect 1564 676 1572 684
rect 1612 676 1620 684
rect 1660 676 1668 684
rect 1772 676 1780 684
rect 1804 676 1812 684
rect 1916 676 1924 684
rect 1980 676 1988 684
rect 2092 676 2100 684
rect 2108 676 2116 684
rect 2220 676 2228 684
rect 2284 676 2292 684
rect 2492 676 2500 684
rect 2556 676 2564 684
rect 2764 676 2772 684
rect 2812 676 2820 684
rect 2876 676 2884 684
rect 3212 676 3220 684
rect 3228 676 3236 684
rect 3340 676 3348 684
rect 3404 676 3412 684
rect 3644 716 3652 724
rect 4028 716 4036 724
rect 4092 716 4100 724
rect 4140 716 4148 724
rect 4236 716 4244 724
rect 4300 716 4308 724
rect 4364 716 4372 724
rect 4428 716 4436 724
rect 4476 716 4484 724
rect 4604 716 4612 724
rect 4716 736 4724 744
rect 5532 756 5540 764
rect 4764 736 4772 744
rect 5484 736 5492 744
rect 5868 736 5876 744
rect 4940 716 4948 724
rect 5388 716 5396 724
rect 5548 716 5556 724
rect 5788 716 5796 724
rect 3516 696 3524 704
rect 3580 696 3588 704
rect 3596 696 3604 704
rect 3724 696 3732 704
rect 3852 696 3860 704
rect 3916 696 3924 704
rect 4012 696 4020 704
rect 4044 696 4052 704
rect 4124 696 4132 704
rect 4204 696 4212 704
rect 4268 696 4276 704
rect 4348 696 4356 704
rect 4380 696 4388 704
rect 4428 696 4436 704
rect 3596 676 3604 684
rect 3676 676 3684 684
rect 3724 676 3732 684
rect 3740 676 3748 684
rect 3788 676 3796 684
rect 3980 676 3988 684
rect 4188 676 4196 684
rect 4236 676 4244 684
rect 4252 676 4260 684
rect 4380 676 4388 684
rect 4492 696 4500 704
rect 4524 696 4532 704
rect 4636 696 4644 704
rect 4684 696 4692 704
rect 4748 696 4756 704
rect 4828 696 4836 704
rect 4844 696 4852 704
rect 4924 696 4932 704
rect 5004 696 5012 704
rect 5036 696 5044 704
rect 5324 696 5332 704
rect 5372 696 5380 704
rect 5580 696 5588 704
rect 5612 696 5620 704
rect 5628 696 5636 704
rect 5740 696 5748 704
rect 5788 696 5796 704
rect 5820 696 5828 704
rect 6172 716 6180 724
rect 5948 696 5956 704
rect 6156 696 6164 704
rect 6252 696 6260 704
rect 4556 676 4564 684
rect 4604 676 4612 684
rect 4636 676 4644 684
rect 4668 676 4676 684
rect 5116 676 5124 684
rect 5148 676 5156 684
rect 5276 676 5284 684
rect 5292 676 5300 684
rect 5468 676 5476 684
rect 5516 676 5524 684
rect 5548 676 5556 684
rect 5564 676 5572 684
rect 5644 676 5652 684
rect 5836 676 5844 684
rect 5916 676 5924 684
rect 5996 676 6004 684
rect 6220 676 6228 684
rect 12 656 20 664
rect 60 656 68 664
rect 124 656 132 664
rect 204 656 212 664
rect 220 656 228 664
rect 300 656 308 664
rect 348 656 356 664
rect 412 656 420 664
rect 428 656 436 664
rect 524 656 532 664
rect 1228 656 1236 664
rect 1452 656 1460 664
rect 2156 656 2164 664
rect 2172 656 2180 664
rect 2268 656 2276 664
rect 2556 656 2564 664
rect 2668 656 2676 664
rect 2860 656 2868 664
rect 3660 656 3668 664
rect 3868 656 3876 664
rect 3980 656 3988 664
rect 4156 656 4164 664
rect 4492 656 4500 664
rect 4716 656 4724 664
rect 4876 656 4884 664
rect 4924 656 4932 664
rect 5292 656 5300 664
rect 5340 656 5348 664
rect 5692 656 5700 664
rect 5708 656 5716 664
rect 5756 656 5764 664
rect 5788 656 5796 664
rect 6060 656 6068 664
rect 6076 656 6084 664
rect 6124 656 6132 664
rect 108 636 116 644
rect 364 636 372 644
rect 508 636 516 644
rect 556 636 564 644
rect 620 636 628 644
rect 668 636 676 644
rect 924 636 932 644
rect 1708 636 1716 644
rect 1884 636 1892 644
rect 1964 636 1972 644
rect 2044 636 2052 644
rect 2380 636 2388 644
rect 2572 636 2580 644
rect 2796 636 2804 644
rect 2972 636 2980 644
rect 3084 636 3092 644
rect 3244 636 3252 644
rect 3292 636 3300 644
rect 3436 636 3444 644
rect 3564 636 3572 644
rect 3756 636 3764 644
rect 3916 636 3924 644
rect 4220 636 4228 644
rect 4300 636 4308 644
rect 4316 636 4324 644
rect 4460 636 4468 644
rect 4572 636 4580 644
rect 4684 636 4692 644
rect 5020 636 5028 644
rect 5228 636 5236 644
rect 5244 636 5252 644
rect 5420 636 5428 644
rect 5580 636 5588 644
rect 3113 606 3121 614
rect 3123 606 3131 614
rect 3133 606 3141 614
rect 3143 606 3151 614
rect 380 576 388 584
rect 796 576 804 584
rect 988 576 996 584
rect 1132 576 1140 584
rect 1260 576 1268 584
rect 2700 576 2708 584
rect 4236 576 4244 584
rect 5052 576 5060 584
rect 5644 576 5652 584
rect 5724 576 5732 584
rect 5884 576 5892 584
rect 6076 576 6084 584
rect 6124 576 6132 584
rect 6204 576 6212 584
rect 6252 576 6260 584
rect 172 556 180 564
rect 348 556 356 564
rect 364 556 372 564
rect 412 556 420 564
rect 476 556 484 564
rect 652 556 660 564
rect 732 556 740 564
rect 1164 556 1172 564
rect 1196 556 1204 564
rect 140 536 148 544
rect 492 536 500 544
rect 556 536 564 544
rect 748 536 756 544
rect 812 536 820 544
rect 1132 536 1140 544
rect 1212 536 1220 544
rect 1324 536 1332 544
rect 1388 536 1396 544
rect 1500 536 1508 544
rect 1516 536 1524 544
rect 1628 556 1636 564
rect 1868 556 1876 564
rect 2060 556 2068 564
rect 2076 556 2084 564
rect 2092 556 2100 564
rect 2268 556 2276 564
rect 2380 556 2388 564
rect 2444 556 2452 564
rect 2652 556 2660 564
rect 2860 556 2868 564
rect 3116 556 3124 564
rect 3340 556 3348 564
rect 3580 556 3588 564
rect 3596 556 3604 564
rect 1676 536 1684 544
rect 1772 536 1780 544
rect 1964 536 1972 544
rect 2108 536 2116 544
rect 2172 536 2180 544
rect 2220 536 2228 544
rect 2252 536 2260 544
rect 2332 536 2340 544
rect 2348 536 2356 544
rect 2380 536 2388 544
rect 2396 536 2404 544
rect 2476 536 2484 544
rect 2492 536 2500 544
rect 2620 536 2628 544
rect 2908 536 2916 544
rect 2956 536 2964 544
rect 3020 536 3028 544
rect 3164 536 3172 544
rect 3180 536 3188 544
rect 3340 536 3348 544
rect 3548 536 3556 544
rect 252 516 260 524
rect 620 516 628 524
rect 700 516 708 524
rect 764 516 772 524
rect 860 516 868 524
rect 924 516 932 524
rect 940 516 948 524
rect 1084 516 1092 524
rect 1148 516 1156 524
rect 1164 516 1172 524
rect 76 500 84 508
rect 588 496 596 504
rect 844 496 852 504
rect 1372 516 1380 524
rect 1404 516 1412 524
rect 1468 516 1476 524
rect 1580 516 1588 524
rect 1724 516 1732 524
rect 1852 516 1860 524
rect 1900 516 1908 524
rect 1948 516 1956 524
rect 1996 516 2004 524
rect 2028 516 2036 524
rect 2124 516 2132 524
rect 1276 496 1284 504
rect 1340 496 1348 504
rect 1452 496 1460 504
rect 1916 496 1924 504
rect 1948 496 1956 504
rect 1980 496 1988 504
rect 2156 496 2164 504
rect 2204 516 2212 524
rect 2236 516 2244 524
rect 2316 516 2324 524
rect 2348 516 2356 524
rect 2492 516 2500 524
rect 2524 516 2532 524
rect 2284 496 2292 504
rect 2620 516 2628 524
rect 2748 516 2756 524
rect 2828 516 2836 524
rect 2892 516 2900 524
rect 2972 516 2980 524
rect 3004 516 3012 524
rect 3036 516 3044 524
rect 3084 516 3092 524
rect 3196 516 3204 524
rect 3260 516 3268 524
rect 3372 516 3380 524
rect 3452 516 3460 524
rect 3500 516 3508 524
rect 2572 496 2580 504
rect 2636 496 2644 504
rect 2780 496 2788 504
rect 2844 496 2852 504
rect 2908 496 2916 504
rect 2924 496 2932 504
rect 3004 496 3012 504
rect 3036 496 3044 504
rect 3068 496 3076 504
rect 3148 496 3156 504
rect 3180 496 3188 504
rect 3356 496 3364 504
rect 908 476 916 484
rect 2012 476 2020 484
rect 2812 476 2820 484
rect 3276 476 3284 484
rect 3388 476 3396 484
rect 3436 476 3444 484
rect 3484 496 3492 504
rect 3596 516 3604 524
rect 3644 556 3652 564
rect 3660 556 3668 564
rect 3676 556 3684 564
rect 3836 556 3844 564
rect 4140 556 4148 564
rect 4172 556 4180 564
rect 4588 556 4596 564
rect 5100 556 5108 564
rect 5228 556 5236 564
rect 5260 556 5268 564
rect 5356 556 5364 564
rect 5372 556 5380 564
rect 5484 556 5492 564
rect 5900 556 5908 564
rect 6140 556 6148 564
rect 3756 536 3764 544
rect 3772 536 3780 544
rect 3852 536 3860 544
rect 3996 536 4004 544
rect 4028 536 4036 544
rect 4060 536 4068 544
rect 4332 536 4340 544
rect 4604 536 4612 544
rect 4652 536 4660 544
rect 4876 536 4884 544
rect 4924 536 4932 544
rect 5212 536 5220 544
rect 5420 536 5428 544
rect 5484 536 5492 544
rect 5548 536 5556 544
rect 5660 536 5668 544
rect 5676 536 5684 544
rect 5740 536 5748 544
rect 5804 536 5812 544
rect 5964 536 5972 544
rect 3676 516 3684 524
rect 3740 516 3748 524
rect 3788 516 3796 524
rect 3916 516 3924 524
rect 4012 516 4020 524
rect 4124 516 4132 524
rect 4140 516 4148 524
rect 4188 516 4196 524
rect 4204 516 4212 524
rect 4252 516 4260 524
rect 4316 516 4324 524
rect 4412 516 4420 524
rect 4460 516 4468 524
rect 4492 516 4500 524
rect 4780 516 4788 524
rect 4812 516 4820 524
rect 4988 516 4996 524
rect 5020 516 5028 524
rect 5068 516 5076 524
rect 5116 516 5124 524
rect 5164 516 5172 524
rect 5212 516 5220 524
rect 3820 496 3828 504
rect 3964 496 3972 504
rect 4060 496 4068 504
rect 4524 496 4532 504
rect 4780 496 4788 504
rect 4828 496 4836 504
rect 4924 496 4932 504
rect 5548 516 5556 524
rect 5580 516 5588 524
rect 5628 516 5636 524
rect 5788 516 5796 524
rect 5852 516 5860 524
rect 5868 516 5876 524
rect 6076 516 6084 524
rect 6284 516 6292 524
rect 5500 496 5508 504
rect 5564 496 5572 504
rect 5724 496 5732 504
rect 5916 496 5924 504
rect 3516 476 3524 484
rect 3932 476 3940 484
rect 4492 476 4500 484
rect 5036 476 5044 484
rect 5596 476 5604 484
rect 5996 476 6004 484
rect 1612 456 1620 464
rect 2044 456 2052 464
rect 3452 456 3460 464
rect 5580 456 5588 464
rect 76 436 84 444
rect 1052 436 1060 444
rect 1372 436 1380 444
rect 1420 436 1428 444
rect 1708 436 1716 444
rect 1740 436 1748 444
rect 1884 436 1892 444
rect 2316 436 2324 444
rect 2524 436 2532 444
rect 2748 436 2756 444
rect 2828 436 2836 444
rect 2972 436 2980 444
rect 3372 436 3380 444
rect 3500 436 3508 444
rect 3612 436 3620 444
rect 3708 436 3716 444
rect 3788 436 3796 444
rect 3916 436 3924 444
rect 4044 436 4052 444
rect 4364 436 4372 444
rect 4428 436 4436 444
rect 4508 436 4516 444
rect 4860 436 4868 444
rect 5068 436 5076 444
rect 5340 436 5348 444
rect 5852 436 5860 444
rect 1577 406 1585 414
rect 1587 406 1595 414
rect 1597 406 1605 414
rect 1607 406 1615 414
rect 4665 406 4673 414
rect 4675 406 4683 414
rect 4685 406 4693 414
rect 4695 406 4703 414
rect 28 376 36 384
rect 284 376 292 384
rect 380 376 388 384
rect 668 376 676 384
rect 732 376 740 384
rect 1836 376 1844 384
rect 2316 376 2324 384
rect 4220 376 4228 384
rect 4524 376 4532 384
rect 5196 376 5204 384
rect 6140 376 6148 384
rect 6172 376 6180 384
rect 988 358 996 366
rect 2460 356 2468 364
rect 1228 336 1236 344
rect 1644 336 1652 344
rect 1788 336 1796 344
rect 1820 336 1828 344
rect 1964 336 1972 344
rect 2636 336 2644 344
rect 2668 336 2676 344
rect 2764 336 2772 344
rect 2796 336 2804 344
rect 2812 336 2820 344
rect 2956 336 2964 344
rect 3532 336 3540 344
rect 4092 356 4100 364
rect 4268 356 4276 364
rect 5372 356 5380 364
rect 5532 356 5540 364
rect 3564 336 3572 344
rect 3612 336 3620 344
rect 3676 336 3684 344
rect 3788 336 3796 344
rect 3932 336 3940 344
rect 4508 336 4516 344
rect 4764 336 4772 344
rect 5276 336 5284 344
rect 5356 336 5364 344
rect 5500 336 5508 344
rect 5644 336 5652 344
rect 5852 336 5860 344
rect 284 312 292 320
rect 668 316 676 324
rect 988 312 996 320
rect 108 296 116 304
rect 316 296 324 304
rect 460 296 468 304
rect 684 296 692 304
rect 812 296 820 304
rect 1308 316 1316 324
rect 1372 316 1380 324
rect 1500 316 1508 324
rect 1564 316 1572 324
rect 1676 316 1684 324
rect 1852 316 1860 324
rect 1868 316 1876 324
rect 1900 316 1908 324
rect 1932 316 1940 324
rect 2156 316 2164 324
rect 2364 316 2372 324
rect 2492 316 2500 324
rect 2540 316 2548 324
rect 2604 316 2612 324
rect 2828 316 2836 324
rect 2988 316 2996 324
rect 3068 316 3076 324
rect 3468 316 3476 324
rect 3532 316 3540 324
rect 3644 316 3652 324
rect 3708 316 3716 324
rect 3820 316 3828 324
rect 3836 316 3844 324
rect 3900 316 3908 324
rect 4428 316 4436 324
rect 4476 316 4484 324
rect 4540 316 4548 324
rect 4684 316 4692 324
rect 4812 316 4820 324
rect 4924 316 4932 324
rect 5004 316 5012 324
rect 5052 316 5060 324
rect 5068 316 5076 324
rect 5324 316 5332 324
rect 5468 316 5476 324
rect 6060 316 6068 324
rect 6092 316 6100 324
rect 6156 316 6164 324
rect 1148 296 1156 304
rect 1276 296 1284 304
rect 1340 296 1348 304
rect 1500 296 1508 304
rect 1564 296 1572 304
rect 1692 296 1700 304
rect 1724 296 1732 304
rect 1756 296 1764 304
rect 1836 296 1844 304
rect 1900 296 1908 304
rect 1948 296 1956 304
rect 1996 296 2004 304
rect 2028 296 2036 304
rect 2236 296 2244 304
rect 2332 296 2340 304
rect 2396 296 2404 304
rect 2556 296 2564 304
rect 2620 296 2628 304
rect 2716 296 2724 304
rect 2764 296 2772 304
rect 220 276 228 284
rect 572 276 580 284
rect 924 276 932 284
rect 1068 276 1076 284
rect 1164 276 1172 284
rect 188 256 196 264
rect 540 256 548 264
rect 892 256 900 264
rect 1260 276 1268 284
rect 1324 276 1332 284
rect 1388 276 1396 284
rect 1404 280 1412 288
rect 1452 276 1460 284
rect 1484 276 1492 284
rect 1516 276 1524 284
rect 1628 276 1636 284
rect 1740 276 1748 284
rect 1916 276 1924 284
rect 2060 276 2068 284
rect 2188 276 2196 284
rect 2252 276 2260 284
rect 2268 276 2276 284
rect 2428 276 2436 284
rect 2508 276 2516 284
rect 2732 276 2740 284
rect 1308 256 1316 264
rect 1612 256 1620 264
rect 1724 256 1732 264
rect 1996 256 2004 264
rect 2028 256 2036 264
rect 2140 256 2148 264
rect 2268 256 2276 264
rect 2428 256 2436 264
rect 2588 256 2596 264
rect 2620 256 2628 264
rect 2668 256 2676 264
rect 2732 256 2740 264
rect 2796 256 2804 264
rect 2844 296 2852 304
rect 2924 296 2932 304
rect 2972 296 2980 304
rect 3004 296 3012 304
rect 3340 296 3348 304
rect 3420 296 3428 304
rect 3468 296 3476 304
rect 3516 296 3524 304
rect 3548 296 3556 304
rect 3660 296 3668 304
rect 3756 296 3764 304
rect 3804 296 3812 304
rect 3868 296 3876 304
rect 3916 296 3924 304
rect 3964 296 3972 304
rect 4028 296 4036 304
rect 4060 296 4068 304
rect 4092 296 4100 304
rect 4172 296 4180 304
rect 4300 296 4308 304
rect 4412 296 4420 304
rect 4492 296 4500 304
rect 4556 296 4564 304
rect 4604 296 4612 304
rect 4668 296 4676 304
rect 4748 296 4756 304
rect 4796 296 4804 304
rect 4908 296 4916 304
rect 5196 296 5204 304
rect 5260 296 5268 304
rect 5340 296 5348 304
rect 5388 296 5396 304
rect 5420 296 5428 304
rect 5484 296 5492 304
rect 5580 296 5588 304
rect 5596 296 5604 304
rect 5612 296 5620 304
rect 5644 296 5652 304
rect 5724 296 5732 304
rect 2924 276 2932 284
rect 3020 276 3028 284
rect 3132 276 3140 284
rect 3196 276 3204 284
rect 3228 276 3236 284
rect 3308 276 3316 284
rect 3420 276 3428 284
rect 3484 276 3492 284
rect 3724 276 3732 284
rect 3756 276 3764 284
rect 3884 276 3892 284
rect 3964 276 3972 284
rect 4044 276 4052 284
rect 4060 274 4068 282
rect 4108 276 4116 284
rect 4156 276 4164 284
rect 4252 276 4260 284
rect 4316 276 4324 284
rect 4332 276 4340 284
rect 4380 276 4388 284
rect 4460 276 4468 284
rect 4620 276 4628 284
rect 4684 276 4692 284
rect 4812 276 4820 284
rect 4844 276 4852 284
rect 4972 276 4980 284
rect 5020 276 5028 284
rect 5100 276 5108 284
rect 5212 276 5220 284
rect 5404 276 5412 284
rect 5436 276 5444 284
rect 5564 276 5572 284
rect 5676 276 5684 284
rect 5708 276 5716 284
rect 5724 276 5732 284
rect 5788 296 5796 304
rect 5852 296 5860 304
rect 5932 296 5940 304
rect 5948 296 5956 304
rect 6012 296 6020 304
rect 6028 296 6036 304
rect 6108 296 6116 304
rect 5788 276 5796 284
rect 5804 276 5812 284
rect 6044 276 6052 284
rect 6108 276 6116 284
rect 2876 256 2884 264
rect 2892 256 2900 264
rect 3052 256 3060 264
rect 3180 256 3188 264
rect 3340 256 3348 264
rect 3516 256 3524 264
rect 3596 256 3604 264
rect 3836 256 3844 264
rect 4140 256 4148 264
rect 4556 256 4564 264
rect 4636 256 4644 264
rect 4876 256 4884 264
rect 5148 256 5156 264
rect 5228 256 5236 264
rect 5260 256 5268 264
rect 5308 256 5316 264
rect 5532 256 5540 264
rect 5772 256 5780 264
rect 5852 256 5860 264
rect 5884 256 5892 264
rect 5900 256 5908 264
rect 6124 256 6132 264
rect 6252 256 6260 264
rect 1084 236 1092 244
rect 1196 236 1204 244
rect 1372 236 1380 244
rect 1436 236 1444 244
rect 1980 236 1988 244
rect 2124 236 2132 244
rect 2156 236 2164 244
rect 2204 236 2212 244
rect 2412 236 2420 244
rect 2540 236 2548 244
rect 2572 236 2580 244
rect 2812 236 2820 244
rect 2940 236 2948 244
rect 3036 236 3044 244
rect 3356 236 3364 244
rect 3660 236 3668 244
rect 3948 236 3956 244
rect 3996 236 4004 244
rect 4348 236 4356 244
rect 4780 236 4788 244
rect 4924 236 4932 244
rect 4988 236 4996 244
rect 5052 236 5060 244
rect 5484 236 5492 244
rect 5644 236 5652 244
rect 5692 236 5700 244
rect 5964 236 5972 244
rect 6236 236 6244 244
rect 3113 206 3121 214
rect 3123 206 3131 214
rect 3133 206 3141 214
rect 3143 206 3151 214
rect 332 176 340 184
rect 764 176 772 184
rect 972 176 980 184
rect 1180 176 1188 184
rect 1356 176 1364 184
rect 1548 176 1556 184
rect 3228 176 3236 184
rect 3564 176 3572 184
rect 3692 176 3700 184
rect 3788 176 3796 184
rect 3980 176 3988 184
rect 4332 176 4340 184
rect 4380 176 4388 184
rect 4460 176 4468 184
rect 4604 176 4612 184
rect 4876 176 4884 184
rect 5020 176 5028 184
rect 5132 176 5140 184
rect 5164 176 5172 184
rect 5500 176 5508 184
rect 5740 176 5748 184
rect 5996 176 6004 184
rect 6156 176 6164 184
rect 6188 176 6196 184
rect 6236 176 6244 184
rect 172 156 180 164
rect 540 156 548 164
rect 988 156 996 164
rect 1084 156 1092 164
rect 1564 156 1572 164
rect 1708 156 1716 164
rect 1756 156 1764 164
rect 1788 156 1796 164
rect 1836 156 1844 164
rect 1980 156 1988 164
rect 2044 156 2052 164
rect 2108 156 2116 164
rect 2204 156 2212 164
rect 2220 156 2228 164
rect 2300 156 2308 164
rect 2332 156 2340 164
rect 2428 156 2436 164
rect 2460 156 2468 164
rect 140 136 148 144
rect 572 136 580 144
rect 780 136 788 144
rect 860 136 868 144
rect 924 136 932 144
rect 1004 136 1012 144
rect 1068 136 1076 144
rect 1132 136 1140 144
rect 1228 136 1236 144
rect 1244 136 1252 144
rect 1276 136 1284 144
rect 1484 136 1492 144
rect 1500 136 1508 144
rect 1612 136 1620 144
rect 1644 136 1652 144
rect 1692 136 1700 144
rect 2316 136 2324 144
rect 2492 136 2500 144
rect 2780 156 2788 164
rect 2972 156 2980 164
rect 3052 156 3060 164
rect 3196 156 3204 164
rect 3244 156 3252 164
rect 3484 156 3492 164
rect 3548 156 3556 164
rect 3964 156 3972 164
rect 4140 156 4148 164
rect 4156 156 4164 164
rect 4284 156 4292 164
rect 4524 156 4532 164
rect 4540 156 4548 164
rect 4620 156 4628 164
rect 4796 156 4804 164
rect 4860 156 4868 164
rect 5036 156 5044 164
rect 5148 156 5156 164
rect 5276 156 5284 164
rect 5372 156 5380 164
rect 5516 156 5524 164
rect 5532 156 5540 164
rect 5756 156 5764 164
rect 6172 156 6180 164
rect 6252 156 6260 164
rect 2652 136 2660 144
rect 252 116 260 124
rect 378 116 386 124
rect 460 116 468 124
rect 876 116 884 124
rect 908 116 916 124
rect 1052 116 1060 124
rect 1116 116 1124 124
rect 76 100 84 108
rect 636 100 644 108
rect 828 96 836 104
rect 908 96 916 104
rect 972 96 980 104
rect 1020 96 1028 104
rect 1164 96 1172 104
rect 1292 116 1300 124
rect 1372 116 1380 124
rect 1404 116 1412 124
rect 1516 116 1524 124
rect 1660 116 1668 124
rect 1804 116 1812 124
rect 1948 116 1956 124
rect 2076 116 2084 124
rect 2140 116 2148 124
rect 2236 116 2244 124
rect 2252 116 2260 124
rect 2268 116 2276 124
rect 2380 116 2388 124
rect 2460 116 2468 124
rect 2492 116 2500 124
rect 2556 116 2564 124
rect 2748 136 2756 144
rect 2860 136 2868 144
rect 2956 136 2964 144
rect 3116 136 3124 144
rect 3196 136 3204 144
rect 3276 136 3284 144
rect 3308 136 3316 144
rect 3468 136 3476 144
rect 3532 136 3540 144
rect 3580 136 3588 144
rect 3676 136 3684 144
rect 3756 132 3764 140
rect 3772 136 3780 144
rect 3820 136 3828 144
rect 3852 136 3860 144
rect 3916 136 3924 144
rect 4124 136 4132 144
rect 4236 136 4244 144
rect 4348 136 4356 144
rect 4444 136 4452 144
rect 4476 136 4484 144
rect 4828 136 4836 144
rect 4972 136 4980 144
rect 5068 136 5076 144
rect 5340 136 5348 144
rect 5388 136 5396 144
rect 5452 136 5460 144
rect 5708 136 5716 144
rect 5932 136 5940 144
rect 6108 136 6116 144
rect 6140 136 6148 144
rect 6220 136 6228 144
rect 1276 96 1284 104
rect 1308 96 1316 104
rect 1324 96 1332 104
rect 1388 96 1396 104
rect 1420 96 1428 104
rect 1452 96 1460 104
rect 1852 96 1860 104
rect 1980 96 1988 104
rect 2060 96 2068 104
rect 2124 96 2132 104
rect 2172 96 2180 104
rect 2284 96 2292 104
rect 2348 96 2356 104
rect 2364 96 2372 104
rect 2476 96 2484 104
rect 2540 96 2548 104
rect 2732 116 2740 124
rect 2812 116 2820 124
rect 3020 116 3028 124
rect 3324 116 3332 124
rect 3388 116 3396 124
rect 3468 116 3476 124
rect 3532 116 3540 124
rect 3644 116 3652 124
rect 3900 116 3908 124
rect 3964 116 3972 124
rect 4044 116 4052 124
rect 4076 116 4084 124
rect 4108 116 4116 124
rect 4124 116 4132 124
rect 4220 116 4228 124
rect 4364 116 4372 124
rect 4412 116 4420 124
rect 4444 116 4452 124
rect 4492 116 4500 124
rect 4524 116 4532 124
rect 4588 116 4596 124
rect 4620 116 4628 124
rect 2796 96 2804 104
rect 2908 96 2916 104
rect 3052 96 3060 104
rect 3372 96 3380 104
rect 3772 96 3780 104
rect 3884 96 3892 104
rect 3948 96 3956 104
rect 4060 96 4068 104
rect 4076 96 4084 104
rect 4220 96 4228 104
rect 4380 96 4388 104
rect 4812 116 4820 124
rect 4860 116 4868 124
rect 4940 116 4948 124
rect 4940 96 4948 104
rect 5068 116 5076 124
rect 5100 116 5108 124
rect 5180 116 5188 124
rect 5228 116 5236 124
rect 5244 116 5252 124
rect 5276 116 5284 124
rect 5132 96 5140 104
rect 5324 116 5332 124
rect 5404 116 5412 124
rect 5468 116 5476 124
rect 5660 116 5668 124
rect 5900 118 5908 126
rect 5964 116 5972 124
rect 5980 116 5988 124
rect 6028 116 6036 124
rect 6060 116 6068 124
rect 6124 116 6132 124
rect 5452 96 5460 104
rect 876 76 884 84
rect 1052 76 1060 84
rect 1132 76 1140 84
rect 1356 76 1364 84
rect 1596 76 1604 84
rect 1884 76 1892 84
rect 1932 76 1940 84
rect 2028 76 2036 84
rect 2092 76 2100 84
rect 2156 76 2164 84
rect 2396 76 2404 84
rect 2508 76 2516 84
rect 2572 76 2580 84
rect 2828 76 2836 84
rect 3004 76 3012 84
rect 3084 76 3092 84
rect 4028 76 4036 84
rect 4492 76 4500 84
rect 4652 76 4660 84
rect 5068 76 5076 84
rect 5548 76 5556 84
rect 5772 76 5780 84
rect 252 54 260 62
rect 2188 56 2196 64
rect 2764 56 2772 64
rect 2924 56 2932 64
rect 5228 56 5236 64
rect 636 36 644 44
rect 2380 36 2388 44
rect 2668 36 2676 44
rect 2876 36 2884 44
rect 2988 36 2996 44
rect 3452 36 3460 44
rect 4748 36 4756 44
rect 5356 36 5364 44
rect 1948 22 1956 30
rect 1577 6 1585 14
rect 1587 6 1595 14
rect 1597 6 1605 14
rect 1607 6 1615 14
rect 4665 6 4673 14
rect 4675 6 4683 14
rect 4685 6 4693 14
rect 4695 6 4703 14
<< metal2 >>
rect 397 4604 403 4643
rect 573 4637 595 4643
rect 141 4577 156 4583
rect 141 4564 147 4577
rect 13 4504 19 4516
rect 93 4504 99 4516
rect 125 4124 131 4136
rect 77 4064 83 4116
rect 173 3984 179 4296
rect 269 4284 275 4536
rect 397 4524 403 4596
rect 573 4563 579 4637
rect 596 4577 611 4583
rect 605 4564 611 4577
rect 573 4557 595 4563
rect 461 4464 467 4536
rect 205 4184 211 4196
rect 301 4183 307 4296
rect 461 4284 467 4456
rect 589 4384 595 4557
rect 637 4504 643 4643
rect 749 4584 755 4643
rect 877 4637 899 4643
rect 669 4544 675 4576
rect 733 4544 739 4576
rect 717 4504 723 4516
rect 733 4304 739 4456
rect 301 4177 380 4183
rect 196 4117 236 4123
rect 205 4084 211 4096
rect 285 3964 291 4116
rect 333 4104 339 4156
rect 349 4104 355 4136
rect 365 4084 371 4116
rect 397 4104 403 4196
rect 477 4164 483 4296
rect 509 4164 515 4276
rect 573 4184 579 4236
rect 653 4164 659 4176
rect 701 4164 707 4296
rect 733 4164 739 4296
rect 429 4144 435 4156
rect 413 4124 419 4136
rect 509 4043 515 4118
rect 493 4037 515 4043
rect 493 3984 499 4037
rect 557 3984 563 4136
rect 269 3904 275 3956
rect 13 3823 19 3856
rect 13 3817 35 3823
rect 29 3644 35 3817
rect 45 3784 51 3856
rect 125 3784 131 3896
rect 173 3884 179 3896
rect 285 3884 291 3896
rect 333 3884 339 3936
rect 244 3877 252 3883
rect 340 3877 355 3883
rect 141 3844 147 3876
rect 157 3784 163 3856
rect 205 3784 211 3876
rect 221 3864 227 3876
rect 317 3844 323 3856
rect 237 3804 243 3836
rect 301 3823 307 3836
rect 285 3817 307 3823
rect 61 3744 67 3756
rect 93 3744 99 3776
rect 253 3763 259 3816
rect 285 3784 291 3817
rect 333 3784 339 3796
rect 244 3757 259 3763
rect 132 3737 140 3743
rect 13 3603 19 3636
rect 45 3604 51 3736
rect 77 3724 83 3736
rect 93 3724 99 3736
rect 125 3604 131 3716
rect 173 3704 179 3716
rect 13 3597 35 3603
rect 29 3544 35 3597
rect 77 3564 83 3596
rect 173 3584 179 3696
rect 205 3604 211 3736
rect 301 3724 307 3776
rect 333 3644 339 3696
rect 205 3564 211 3596
rect 349 3564 355 3877
rect 365 3844 371 3876
rect 381 3844 387 3916
rect 445 3744 451 3916
rect 461 3884 467 3916
rect 525 3904 531 3916
rect 509 3864 515 3876
rect 461 3784 467 3796
rect 420 3737 435 3743
rect 429 3723 435 3737
rect 468 3737 476 3743
rect 509 3724 515 3836
rect 525 3764 531 3896
rect 605 3884 611 4096
rect 637 4084 643 4096
rect 781 4004 787 4516
rect 845 4464 851 4536
rect 893 4384 899 4637
rect 980 4577 995 4583
rect 989 4564 995 4577
rect 973 4384 979 4556
rect 1021 4544 1027 4576
rect 1053 4504 1059 4643
rect 1165 4637 1187 4643
rect 1149 4577 1164 4583
rect 1069 4544 1075 4576
rect 1149 4564 1155 4577
rect 1181 4563 1187 4637
rect 1373 4577 1388 4583
rect 1373 4564 1379 4577
rect 1165 4557 1187 4563
rect 1085 4504 1091 4516
rect 1117 4484 1123 4496
rect 941 4324 947 4336
rect 1005 4304 1011 4316
rect 1085 4304 1091 4436
rect 1165 4384 1171 4557
rect 1261 4524 1267 4556
rect 1277 4464 1283 4536
rect 813 4224 819 4236
rect 861 4204 867 4276
rect 868 4177 883 4183
rect 877 4164 883 4177
rect 877 4024 883 4076
rect 909 4064 915 4116
rect 925 4084 931 4296
rect 1085 4284 1091 4296
rect 1069 4264 1075 4276
rect 973 4144 979 4156
rect 957 4104 963 4136
rect 989 4124 995 4256
rect 1037 4217 1091 4223
rect 1037 4163 1043 4217
rect 1021 4157 1043 4163
rect 1021 4144 1027 4157
rect 1037 4124 1043 4136
rect 1053 4124 1059 4196
rect 1085 4124 1091 4217
rect 1101 4184 1107 4216
rect 973 4064 979 4116
rect 685 3904 691 3916
rect 589 3744 595 3776
rect 429 3717 444 3723
rect 397 3703 403 3716
rect 589 3704 595 3716
rect 397 3697 412 3703
rect 77 3524 83 3556
rect 141 3464 147 3476
rect 205 3444 211 3480
rect 285 3483 291 3536
rect 397 3484 403 3496
rect 413 3484 419 3516
rect 429 3504 435 3636
rect 493 3584 499 3596
rect 493 3484 499 3496
rect 285 3477 332 3483
rect 221 3464 227 3476
rect 349 3464 355 3476
rect 61 2984 67 3318
rect 77 3084 83 3336
rect 125 3324 131 3376
rect 173 3324 179 3436
rect 189 3364 195 3376
rect 205 3164 211 3336
rect 221 3283 227 3456
rect 269 3324 275 3436
rect 333 3404 339 3436
rect 429 3384 435 3476
rect 525 3443 531 3516
rect 541 3484 547 3696
rect 605 3683 611 3876
rect 813 3864 819 3936
rect 637 3784 643 3816
rect 669 3744 675 3856
rect 813 3804 819 3856
rect 701 3726 707 3796
rect 829 3744 835 3776
rect 877 3744 883 4016
rect 893 3944 899 4036
rect 701 3717 707 3718
rect 589 3677 611 3683
rect 557 3544 563 3676
rect 557 3524 563 3536
rect 573 3484 579 3496
rect 525 3437 547 3443
rect 365 3324 371 3376
rect 429 3344 435 3376
rect 461 3303 467 3436
rect 541 3404 547 3437
rect 509 3344 515 3356
rect 461 3297 483 3303
rect 221 3277 243 3283
rect 93 3104 99 3116
rect 205 3064 211 3076
rect 237 2984 243 3277
rect 445 3224 451 3236
rect 349 3184 355 3216
rect 413 3184 419 3196
rect 365 3144 371 3156
rect 317 3104 323 3136
rect 413 3124 419 3156
rect 333 3083 339 3116
rect 349 3104 355 3116
rect 420 3097 435 3103
rect 317 3077 339 3083
rect 269 3023 275 3076
rect 285 3044 291 3056
rect 253 3017 275 3023
rect 253 2984 259 3017
rect 13 2904 19 2936
rect 29 2924 35 2956
rect 84 2937 99 2943
rect 93 2924 99 2937
rect 13 2544 19 2896
rect 77 2704 83 2856
rect 125 2784 131 2916
rect 141 2864 147 2936
rect 189 2864 195 2916
rect 221 2904 227 2936
rect 301 2924 307 3036
rect 317 2904 323 3077
rect 429 2984 435 3097
rect 221 2784 227 2876
rect 253 2864 259 2876
rect 317 2844 323 2896
rect 333 2823 339 2936
rect 477 2923 483 3297
rect 525 3244 531 3256
rect 525 3104 531 3236
rect 541 3204 547 3336
rect 557 3163 563 3336
rect 541 3157 563 3163
rect 493 2924 499 3036
rect 509 2944 515 3016
rect 468 2917 483 2923
rect 500 2917 508 2923
rect 397 2904 403 2916
rect 333 2817 355 2823
rect 93 2684 99 2736
rect 141 2664 147 2776
rect 93 2584 99 2636
rect 157 2584 163 2716
rect 221 2684 227 2696
rect 237 2684 243 2756
rect 292 2717 307 2723
rect 93 2563 99 2576
rect 84 2557 99 2563
rect 173 2563 179 2676
rect 173 2557 195 2563
rect 141 2544 147 2556
rect 20 2517 28 2523
rect 13 2304 19 2516
rect 45 2384 51 2536
rect 141 2384 147 2536
rect 189 2524 195 2557
rect 237 2543 243 2676
rect 269 2664 275 2696
rect 285 2624 291 2636
rect 253 2564 259 2616
rect 301 2604 307 2717
rect 349 2723 355 2817
rect 349 2717 387 2723
rect 333 2704 339 2716
rect 365 2704 371 2717
rect 381 2704 387 2717
rect 333 2584 339 2676
rect 349 2604 355 2696
rect 397 2684 403 2856
rect 413 2764 419 2896
rect 484 2877 499 2883
rect 493 2863 499 2877
rect 493 2857 515 2863
rect 509 2844 515 2857
rect 525 2844 531 3076
rect 541 3004 547 3157
rect 557 3124 563 3136
rect 573 3124 579 3456
rect 589 3344 595 3677
rect 605 3524 611 3616
rect 621 3584 627 3636
rect 637 3504 643 3576
rect 653 3484 659 3596
rect 669 3504 675 3696
rect 749 3584 755 3596
rect 765 3563 771 3596
rect 733 3557 771 3563
rect 589 3304 595 3336
rect 605 3324 611 3476
rect 621 3464 627 3476
rect 669 3463 675 3496
rect 701 3484 707 3516
rect 733 3464 739 3557
rect 797 3524 803 3536
rect 813 3504 819 3716
rect 861 3544 867 3736
rect 877 3584 883 3596
rect 893 3544 899 3936
rect 909 3924 915 4056
rect 989 4044 995 4076
rect 909 3904 915 3916
rect 941 3884 947 3996
rect 1005 3904 1011 4116
rect 1021 4084 1027 4096
rect 1085 4064 1091 4096
rect 1101 4084 1107 4156
rect 1117 4044 1123 4256
rect 1149 4064 1155 4116
rect 1021 3904 1027 3916
rect 909 3784 915 3836
rect 925 3744 931 3756
rect 973 3743 979 3836
rect 973 3737 988 3743
rect 909 3664 915 3696
rect 941 3684 947 3696
rect 957 3564 963 3736
rect 989 3703 995 3716
rect 989 3697 1011 3703
rect 1005 3684 1011 3697
rect 973 3644 979 3656
rect 781 3484 787 3496
rect 669 3457 691 3463
rect 621 3404 627 3456
rect 653 3443 659 3456
rect 685 3443 691 3457
rect 653 3437 675 3443
rect 685 3437 716 3443
rect 669 3423 675 3437
rect 797 3443 803 3476
rect 781 3437 803 3443
rect 781 3423 787 3437
rect 669 3417 787 3423
rect 685 3344 691 3376
rect 685 3324 691 3336
rect 781 3304 787 3336
rect 717 3244 723 3296
rect 749 3284 755 3296
rect 589 3184 595 3196
rect 589 3124 595 3176
rect 605 3084 611 3156
rect 621 3084 627 3096
rect 685 3084 691 3236
rect 557 3044 563 3056
rect 557 2964 563 3036
rect 493 2703 499 2836
rect 525 2703 531 2756
rect 541 2724 547 2916
rect 557 2764 563 2936
rect 573 2924 579 3076
rect 637 3044 643 3076
rect 685 3064 691 3076
rect 701 3064 707 3096
rect 717 3084 723 3116
rect 589 2917 604 2923
rect 589 2864 595 2917
rect 573 2723 579 2796
rect 564 2717 579 2723
rect 477 2697 499 2703
rect 509 2697 531 2703
rect 372 2677 380 2683
rect 228 2537 243 2543
rect 317 2524 323 2576
rect 333 2324 339 2536
rect 141 2264 147 2296
rect 301 2284 307 2316
rect 349 2304 355 2336
rect 269 2263 275 2276
rect 253 2257 275 2263
rect 253 2244 259 2257
rect 301 2164 307 2276
rect 333 2264 339 2276
rect 365 2204 371 2536
rect 429 2524 435 2636
rect 381 2284 387 2296
rect 413 2264 419 2356
rect 445 2283 451 2616
rect 477 2603 483 2697
rect 509 2684 515 2697
rect 493 2644 499 2676
rect 509 2624 515 2636
rect 461 2597 483 2603
rect 461 2564 467 2597
rect 509 2584 515 2616
rect 461 2524 467 2536
rect 477 2323 483 2396
rect 493 2323 499 2556
rect 477 2317 499 2323
rect 477 2304 483 2317
rect 445 2277 467 2283
rect 429 2244 435 2256
rect 397 2184 403 2216
rect 13 1984 19 1996
rect 77 1784 83 2096
rect 109 1724 115 1896
rect 125 1884 131 2136
rect 141 2126 147 2156
rect 253 2144 259 2156
rect 141 2117 147 2118
rect 141 1902 147 1916
rect 221 1864 227 1876
rect 173 1744 179 1856
rect 237 1843 243 1896
rect 253 1844 259 1856
rect 221 1837 243 1843
rect 173 1724 179 1736
rect 109 1704 115 1716
rect 189 1704 195 1836
rect 221 1784 227 1837
rect 237 1744 243 1756
rect 157 1684 163 1696
rect 173 1664 179 1696
rect 13 1384 19 1516
rect 45 1504 51 1516
rect 61 1384 67 1476
rect 93 1464 99 1536
rect 205 1384 211 1476
rect 237 1384 243 1736
rect 269 1544 275 2116
rect 301 2104 307 2116
rect 317 2104 323 2116
rect 349 2104 355 2156
rect 429 2144 435 2156
rect 388 2137 403 2143
rect 397 2124 403 2137
rect 461 2143 467 2277
rect 509 2264 515 2356
rect 525 2344 531 2676
rect 541 2584 547 2716
rect 573 2664 579 2696
rect 589 2643 595 2716
rect 605 2664 611 2836
rect 564 2637 595 2643
rect 621 2624 627 3016
rect 653 2944 659 2956
rect 669 2924 675 3036
rect 733 2964 739 3156
rect 765 3123 771 3236
rect 797 3144 803 3236
rect 813 3123 819 3496
rect 861 3484 867 3536
rect 893 3504 899 3516
rect 829 3464 835 3476
rect 868 3457 883 3463
rect 829 3343 835 3356
rect 829 3337 851 3343
rect 845 3324 851 3337
rect 877 3264 883 3457
rect 893 3384 899 3476
rect 909 3384 915 3536
rect 989 3524 995 3676
rect 1021 3583 1027 3896
rect 1037 3884 1043 3976
rect 1069 3884 1075 3956
rect 1085 3917 1100 3923
rect 1085 3904 1091 3917
rect 1069 3864 1075 3876
rect 1085 3864 1091 3876
rect 1117 3843 1123 3976
rect 1133 3924 1139 3976
rect 1149 3904 1155 3916
rect 1165 3903 1171 4036
rect 1197 4024 1203 4296
rect 1245 4284 1251 4456
rect 1261 4224 1267 4296
rect 1277 4123 1283 4276
rect 1261 4117 1283 4123
rect 1261 4104 1267 4117
rect 1293 4104 1299 4236
rect 1325 4164 1331 4236
rect 1341 4184 1347 4476
rect 1405 4384 1411 4643
rect 1629 4624 1635 4643
rect 1709 4624 1715 4643
rect 1757 4624 1763 4643
rect 1837 4637 1859 4643
rect 1421 4384 1427 4496
rect 1501 4464 1507 4536
rect 1549 4384 1555 4616
rect 1725 4584 1731 4616
rect 1789 4557 1804 4563
rect 1789 4544 1795 4557
rect 1597 4504 1603 4536
rect 1613 4444 1619 4536
rect 1700 4517 1715 4523
rect 1629 4504 1635 4516
rect 1645 4504 1651 4516
rect 1677 4504 1683 4516
rect 1576 4406 1577 4414
rect 1585 4406 1587 4414
rect 1595 4406 1597 4414
rect 1605 4406 1607 4414
rect 1615 4406 1624 4414
rect 1533 4363 1539 4376
rect 1533 4357 1571 4363
rect 1380 4297 1395 4303
rect 1373 4184 1379 4276
rect 1389 4144 1395 4297
rect 1485 4284 1491 4336
rect 1501 4284 1507 4296
rect 1405 4184 1411 4256
rect 1469 4184 1475 4216
rect 1332 4137 1347 4143
rect 1341 4124 1347 4137
rect 1309 4104 1315 4116
rect 1389 4064 1395 4136
rect 1341 4024 1347 4036
rect 1181 3924 1187 3976
rect 1229 3937 1276 3943
rect 1229 3924 1235 3937
rect 1252 3917 1260 3923
rect 1165 3897 1219 3903
rect 1133 3864 1139 3896
rect 1213 3884 1219 3897
rect 1117 3837 1139 3843
rect 1037 3644 1043 3756
rect 1053 3744 1059 3836
rect 1117 3764 1123 3776
rect 1085 3744 1091 3756
rect 1069 3724 1075 3736
rect 1101 3723 1107 3756
rect 1133 3744 1139 3837
rect 1149 3744 1155 3876
rect 1293 3863 1299 3996
rect 1357 3984 1363 4056
rect 1453 4024 1459 4156
rect 1485 4083 1491 4256
rect 1549 4224 1555 4296
rect 1565 4283 1571 4357
rect 1645 4323 1651 4436
rect 1661 4364 1667 4476
rect 1677 4384 1683 4476
rect 1629 4317 1651 4323
rect 1565 4277 1603 4283
rect 1501 4124 1507 4136
rect 1469 4077 1491 4083
rect 1389 3924 1395 3996
rect 1405 3884 1411 3936
rect 1437 3903 1443 3996
rect 1453 3924 1459 3996
rect 1437 3897 1459 3903
rect 1357 3863 1363 3876
rect 1293 3857 1315 3863
rect 1197 3844 1203 3856
rect 1165 3784 1171 3836
rect 1181 3743 1187 3836
rect 1261 3764 1267 3856
rect 1245 3757 1260 3763
rect 1181 3737 1212 3743
rect 1085 3717 1107 3723
rect 1037 3624 1043 3636
rect 1053 3624 1059 3696
rect 1021 3577 1043 3583
rect 925 3424 931 3516
rect 973 3504 979 3516
rect 1005 3463 1011 3536
rect 1037 3504 1043 3577
rect 1069 3563 1075 3696
rect 1085 3604 1091 3717
rect 1101 3684 1107 3696
rect 1060 3557 1075 3563
rect 1021 3484 1027 3496
rect 1085 3483 1091 3576
rect 1101 3484 1107 3676
rect 1117 3564 1123 3696
rect 1133 3584 1139 3736
rect 1149 3524 1155 3716
rect 1213 3703 1219 3716
rect 1245 3704 1251 3757
rect 1277 3744 1283 3776
rect 1309 3744 1315 3857
rect 1341 3857 1363 3863
rect 1341 3844 1347 3857
rect 1437 3844 1443 3876
rect 1453 3844 1459 3897
rect 1469 3764 1475 4077
rect 1517 4024 1523 4136
rect 1565 4123 1571 4277
rect 1597 4264 1603 4277
rect 1581 4143 1587 4256
rect 1629 4184 1635 4317
rect 1693 4303 1699 4416
rect 1652 4297 1699 4303
rect 1693 4184 1699 4236
rect 1709 4184 1715 4517
rect 1805 4523 1811 4536
rect 1796 4517 1811 4523
rect 1757 4183 1763 4356
rect 1773 4304 1779 4356
rect 1789 4324 1795 4496
rect 1757 4177 1779 4183
rect 1613 4143 1619 4156
rect 1581 4137 1619 4143
rect 1565 4117 1580 4123
rect 1597 4083 1603 4116
rect 1533 4077 1603 4083
rect 1533 4064 1539 4077
rect 1485 3937 1539 3943
rect 1485 3904 1491 3937
rect 1533 3924 1539 3937
rect 1549 3904 1555 4056
rect 1629 4043 1635 4176
rect 1677 4124 1683 4156
rect 1741 4144 1747 4156
rect 1652 4117 1667 4123
rect 1629 4037 1651 4043
rect 1576 4006 1577 4014
rect 1585 4006 1587 4014
rect 1595 4006 1597 4014
rect 1605 4006 1607 4014
rect 1615 4006 1624 4014
rect 1485 3784 1491 3856
rect 1309 3717 1324 3723
rect 1213 3697 1235 3703
rect 1165 3684 1171 3696
rect 1229 3684 1235 3697
rect 1181 3624 1187 3676
rect 1197 3544 1203 3556
rect 1117 3504 1123 3516
rect 1076 3477 1091 3483
rect 1117 3483 1123 3496
rect 1165 3483 1171 3516
rect 1181 3504 1187 3516
rect 1117 3477 1139 3483
rect 1165 3477 1187 3483
rect 1005 3457 1020 3463
rect 957 3344 963 3396
rect 989 3324 995 3436
rect 1037 3424 1043 3476
rect 973 3304 979 3316
rect 877 3204 883 3236
rect 765 3117 787 3123
rect 765 3064 771 3096
rect 781 2964 787 3117
rect 797 3117 819 3123
rect 797 3083 803 3117
rect 797 3077 819 3083
rect 813 2964 819 3077
rect 813 2944 819 2956
rect 829 2944 835 3116
rect 845 3084 851 3196
rect 877 3124 883 3196
rect 1005 3144 1011 3416
rect 1069 3404 1075 3476
rect 1133 3464 1139 3477
rect 1181 3464 1187 3477
rect 1213 3483 1219 3576
rect 1229 3504 1235 3536
rect 1261 3504 1267 3696
rect 1309 3643 1315 3717
rect 1293 3637 1315 3643
rect 1293 3524 1299 3637
rect 1277 3504 1283 3516
rect 1293 3484 1299 3496
rect 1309 3484 1315 3536
rect 1213 3477 1228 3483
rect 1197 3463 1203 3476
rect 1197 3457 1219 3463
rect 1117 3404 1123 3456
rect 1149 3443 1155 3456
rect 1133 3437 1171 3443
rect 989 3124 995 3136
rect 909 3084 915 3116
rect 941 3084 947 3116
rect 717 2884 723 2896
rect 669 2784 675 2836
rect 637 2704 643 2716
rect 669 2704 675 2756
rect 749 2702 755 2716
rect 653 2664 659 2676
rect 685 2624 691 2676
rect 525 2324 531 2336
rect 541 2324 547 2476
rect 541 2284 547 2316
rect 557 2304 563 2556
rect 573 2304 579 2516
rect 461 2137 483 2143
rect 372 2117 387 2123
rect 381 2003 387 2117
rect 429 2064 435 2116
rect 477 2103 483 2137
rect 557 2104 563 2276
rect 573 2264 579 2276
rect 573 2104 579 2116
rect 461 2097 483 2103
rect 397 2003 403 2016
rect 381 1997 403 2003
rect 349 1904 355 1976
rect 397 1924 403 1997
rect 413 1924 419 1996
rect 429 1904 435 1916
rect 372 1897 380 1903
rect 349 1884 355 1896
rect 333 1764 339 1876
rect 365 1724 371 1876
rect 461 1863 467 2097
rect 605 2064 611 2576
rect 621 2564 627 2616
rect 749 2564 755 2656
rect 804 2537 819 2543
rect 621 2364 627 2516
rect 637 2404 643 2536
rect 637 2324 643 2396
rect 653 2344 659 2456
rect 669 2424 675 2516
rect 717 2504 723 2516
rect 653 2284 659 2336
rect 669 2284 675 2356
rect 717 2324 723 2496
rect 749 2364 755 2516
rect 781 2504 787 2516
rect 765 2444 771 2496
rect 765 2384 771 2416
rect 733 2304 739 2316
rect 749 2284 755 2356
rect 685 2184 691 2216
rect 701 2144 707 2236
rect 724 2117 739 2123
rect 733 2104 739 2117
rect 765 2104 771 2376
rect 781 2284 787 2296
rect 797 2284 803 2396
rect 813 2384 819 2537
rect 829 2424 835 2556
rect 845 2544 851 2916
rect 861 2684 867 3076
rect 925 3064 931 3080
rect 957 3064 963 3116
rect 1021 3104 1027 3396
rect 1037 3324 1043 3376
rect 1069 3343 1075 3356
rect 1069 3337 1091 3343
rect 1085 3324 1091 3337
rect 980 3097 988 3103
rect 925 3037 963 3043
rect 877 2943 883 3016
rect 893 2963 899 3036
rect 925 3024 931 3037
rect 893 2957 915 2963
rect 877 2937 892 2943
rect 877 2904 883 2916
rect 893 2824 899 2936
rect 909 2903 915 2957
rect 941 2924 947 3016
rect 957 2943 963 3037
rect 973 3024 979 3096
rect 957 2937 972 2943
rect 909 2897 931 2903
rect 925 2884 931 2897
rect 957 2824 963 2876
rect 973 2864 979 2916
rect 1005 2883 1011 3016
rect 1037 2983 1043 3316
rect 1053 3304 1059 3316
rect 1069 3284 1075 3316
rect 1101 3284 1107 3396
rect 1133 3343 1139 3437
rect 1165 3364 1171 3437
rect 1181 3344 1187 3396
rect 1213 3363 1219 3457
rect 1261 3384 1267 3396
rect 1236 3377 1244 3383
rect 1309 3383 1315 3476
rect 1325 3424 1331 3696
rect 1341 3524 1347 3596
rect 1357 3483 1363 3556
rect 1373 3544 1379 3736
rect 1389 3724 1395 3736
rect 1405 3704 1411 3716
rect 1421 3524 1427 3736
rect 1437 3564 1443 3756
rect 1485 3724 1491 3736
rect 1469 3544 1475 3596
rect 1485 3584 1491 3676
rect 1437 3517 1468 3523
rect 1405 3504 1411 3516
rect 1437 3503 1443 3517
rect 1428 3497 1443 3503
rect 1460 3497 1475 3503
rect 1373 3484 1379 3496
rect 1341 3477 1363 3483
rect 1341 3464 1347 3477
rect 1309 3377 1331 3383
rect 1213 3357 1235 3363
rect 1117 3337 1139 3343
rect 1117 3324 1123 3337
rect 1085 3244 1091 3276
rect 1133 3244 1139 3316
rect 1069 3184 1075 3236
rect 1069 3137 1100 3143
rect 1069 3124 1075 3137
rect 1021 2977 1043 2983
rect 1021 2924 1027 2977
rect 1053 2964 1059 3076
rect 1085 3024 1091 3076
rect 1117 3024 1123 3196
rect 1149 3184 1155 3336
rect 1165 3304 1171 3316
rect 1149 3124 1155 3176
rect 1181 3124 1187 3296
rect 1197 3224 1203 3316
rect 1229 3304 1235 3357
rect 1245 3344 1251 3356
rect 1277 3344 1283 3376
rect 1293 3304 1299 3316
rect 1229 3183 1235 3296
rect 1252 3197 1267 3203
rect 1213 3177 1235 3183
rect 1197 3144 1203 3156
rect 1213 3103 1219 3177
rect 1261 3163 1267 3197
rect 1309 3184 1315 3356
rect 1325 3183 1331 3377
rect 1357 3304 1363 3456
rect 1373 3303 1379 3456
rect 1389 3357 1420 3363
rect 1389 3324 1395 3357
rect 1421 3304 1427 3316
rect 1373 3297 1388 3303
rect 1348 3277 1372 3283
rect 1325 3177 1347 3183
rect 1261 3157 1283 3163
rect 1229 3124 1235 3156
rect 1245 3144 1251 3156
rect 1261 3124 1267 3136
rect 1277 3104 1283 3157
rect 1213 3097 1235 3103
rect 1149 3084 1155 3096
rect 1069 2957 1084 2963
rect 1037 2924 1043 2936
rect 1069 2924 1075 2957
rect 1117 2944 1123 2956
rect 1085 2924 1091 2936
rect 1133 2904 1139 3036
rect 1149 2944 1155 2956
rect 1037 2883 1043 2896
rect 1005 2877 1043 2883
rect 893 2764 899 2776
rect 877 2724 883 2736
rect 909 2684 915 2716
rect 925 2624 931 2816
rect 973 2804 979 2856
rect 957 2744 963 2756
rect 1069 2743 1075 2796
rect 1101 2784 1107 2836
rect 1117 2824 1123 2836
rect 1069 2737 1084 2743
rect 1117 2724 1123 2736
rect 1005 2704 1011 2716
rect 1133 2704 1139 2856
rect 1149 2824 1155 2936
rect 1165 2924 1171 3096
rect 1181 3044 1187 3096
rect 1181 2884 1187 2916
rect 1044 2677 1052 2683
rect 941 2544 947 2556
rect 989 2544 995 2596
rect 845 2384 851 2516
rect 877 2464 883 2496
rect 893 2464 899 2536
rect 973 2526 979 2536
rect 973 2517 979 2518
rect 909 2424 915 2516
rect 845 2357 883 2363
rect 829 2324 835 2356
rect 845 2324 851 2357
rect 877 2343 883 2357
rect 877 2337 915 2343
rect 861 2324 867 2336
rect 893 2304 899 2316
rect 909 2304 915 2337
rect 820 2297 844 2303
rect 925 2264 931 2356
rect 941 2344 947 2416
rect 989 2304 995 2476
rect 1021 2283 1027 2496
rect 1069 2484 1075 2676
rect 1101 2584 1107 2696
rect 1165 2683 1171 2836
rect 1181 2744 1187 2816
rect 1197 2723 1203 3076
rect 1213 2944 1219 2976
rect 1229 2944 1235 3097
rect 1309 3064 1315 3076
rect 1309 2944 1315 2956
rect 1341 2944 1347 3177
rect 1357 3104 1363 3216
rect 1389 3104 1395 3256
rect 1357 2924 1363 3036
rect 1389 3024 1395 3096
rect 1252 2917 1260 2923
rect 1229 2897 1244 2903
rect 1229 2784 1235 2897
rect 1316 2877 1331 2883
rect 1213 2744 1219 2756
rect 1188 2717 1203 2723
rect 1229 2704 1235 2716
rect 1245 2684 1251 2716
rect 1149 2677 1171 2683
rect 1133 2624 1139 2676
rect 1117 2564 1123 2576
rect 1149 2544 1155 2677
rect 1261 2664 1267 2836
rect 1277 2664 1283 2876
rect 1325 2804 1331 2877
rect 1309 2704 1315 2776
rect 1165 2524 1171 2536
rect 1149 2504 1155 2516
rect 1021 2277 1043 2283
rect 804 2257 819 2263
rect 797 2224 803 2236
rect 813 2224 819 2257
rect 797 2144 803 2216
rect 813 2164 819 2196
rect 765 2064 771 2096
rect 477 2037 515 2043
rect 477 2024 483 2037
rect 509 2024 515 2037
rect 477 1884 483 1996
rect 493 1984 499 2016
rect 541 1924 547 1976
rect 461 1857 483 1863
rect 477 1804 483 1857
rect 509 1764 515 1876
rect 557 1843 563 2056
rect 621 1963 627 1976
rect 621 1957 643 1963
rect 589 1904 595 1916
rect 557 1837 579 1843
rect 477 1744 483 1756
rect 541 1723 547 1836
rect 557 1764 563 1816
rect 532 1717 547 1723
rect 301 1524 307 1636
rect 365 1584 371 1716
rect 493 1704 499 1716
rect 429 1584 435 1696
rect 301 1484 307 1516
rect 317 1384 323 1416
rect 61 1344 67 1376
rect 189 1344 195 1356
rect 13 1304 19 1316
rect 45 1184 51 1336
rect 317 1324 323 1336
rect 285 1317 300 1323
rect 125 1184 131 1316
rect 157 1184 163 1216
rect 285 1184 291 1317
rect 365 1284 371 1536
rect 397 1504 403 1516
rect 525 1504 531 1616
rect 541 1524 547 1536
rect 573 1524 579 1837
rect 589 1744 595 1836
rect 605 1784 611 1896
rect 621 1844 627 1856
rect 637 1844 643 1957
rect 653 1824 659 1916
rect 669 1903 675 1976
rect 781 1944 787 2016
rect 733 1924 739 1936
rect 829 1924 835 2036
rect 845 2024 851 2116
rect 733 1917 736 1924
rect 669 1897 684 1903
rect 669 1844 675 1876
rect 701 1824 707 1876
rect 621 1784 627 1796
rect 637 1743 643 1796
rect 685 1784 691 1816
rect 717 1804 723 1916
rect 845 1884 851 1896
rect 765 1864 771 1876
rect 628 1737 643 1743
rect 669 1724 675 1756
rect 717 1744 723 1756
rect 765 1744 771 1856
rect 861 1784 867 2116
rect 893 2104 899 2256
rect 1037 2224 1043 2277
rect 1085 2184 1091 2196
rect 893 1904 899 2016
rect 909 1984 915 2136
rect 925 2124 931 2136
rect 957 2063 963 2076
rect 941 2057 963 2063
rect 941 2024 947 2057
rect 973 2004 979 2096
rect 1021 2084 1027 2136
rect 1101 2123 1107 2496
rect 1149 2144 1155 2476
rect 1181 2383 1187 2576
rect 1229 2564 1235 2656
rect 1213 2524 1219 2556
rect 1245 2504 1251 2656
rect 1293 2584 1299 2656
rect 1309 2564 1315 2696
rect 1341 2683 1347 2896
rect 1373 2703 1379 2936
rect 1389 2704 1395 2776
rect 1364 2697 1379 2703
rect 1389 2684 1395 2696
rect 1405 2684 1411 3276
rect 1421 3264 1427 3296
rect 1437 3264 1443 3396
rect 1469 3363 1475 3497
rect 1485 3384 1491 3496
rect 1501 3404 1507 3816
rect 1517 3764 1523 3876
rect 1565 3784 1571 3856
rect 1517 3503 1523 3716
rect 1533 3524 1539 3616
rect 1549 3544 1555 3716
rect 1581 3664 1587 3876
rect 1597 3684 1603 3896
rect 1645 3884 1651 4037
rect 1661 4024 1667 4117
rect 1693 4064 1699 4136
rect 1741 4043 1747 4096
rect 1757 4064 1763 4156
rect 1773 4144 1779 4177
rect 1773 4084 1779 4136
rect 1789 4124 1795 4316
rect 1805 4244 1811 4517
rect 1821 4284 1827 4336
rect 1853 4223 1859 4637
rect 1901 4584 1907 4643
rect 1949 4637 1971 4643
rect 1949 4584 1955 4616
rect 1965 4584 1971 4637
rect 1997 4624 2003 4643
rect 2013 4637 2035 4643
rect 2013 4584 2019 4637
rect 2093 4584 2099 4643
rect 1997 4444 2003 4516
rect 2045 4504 2051 4516
rect 1901 4283 1907 4356
rect 1933 4304 1939 4356
rect 1901 4277 1916 4283
rect 1981 4264 1987 4296
rect 1997 4284 2003 4296
rect 1837 4217 1859 4223
rect 1837 4184 1843 4217
rect 1885 4184 1891 4256
rect 1805 4117 1843 4123
rect 1805 4103 1811 4117
rect 1789 4097 1811 4103
rect 1789 4063 1795 4097
rect 1821 4064 1827 4096
rect 1773 4057 1795 4063
rect 1773 4043 1779 4057
rect 1741 4037 1779 4043
rect 1693 3984 1699 4036
rect 1725 3997 1795 4003
rect 1613 3744 1619 3836
rect 1693 3763 1699 3916
rect 1725 3904 1731 3997
rect 1757 3923 1763 3976
rect 1789 3943 1795 3997
rect 1805 3984 1811 4056
rect 1837 4044 1843 4117
rect 1869 4104 1875 4116
rect 1885 4064 1891 4116
rect 1901 4064 1907 4256
rect 2029 4177 2044 4183
rect 1780 3937 1795 3943
rect 1757 3917 1779 3923
rect 1773 3883 1779 3917
rect 1821 3904 1827 4036
rect 1853 3963 1859 4056
rect 1853 3957 1907 3963
rect 1773 3877 1795 3883
rect 1789 3863 1795 3877
rect 1789 3857 1811 3863
rect 1709 3784 1715 3836
rect 1741 3823 1747 3836
rect 1773 3823 1779 3856
rect 1741 3817 1779 3823
rect 1693 3757 1715 3763
rect 1661 3724 1667 3756
rect 1613 3664 1619 3696
rect 1576 3606 1577 3614
rect 1585 3606 1587 3614
rect 1595 3606 1597 3614
rect 1605 3606 1607 3614
rect 1615 3606 1624 3614
rect 1597 3524 1603 3536
rect 1517 3497 1532 3503
rect 1517 3384 1523 3456
rect 1533 3364 1539 3456
rect 1469 3357 1491 3363
rect 1437 2924 1443 3016
rect 1421 2684 1427 2856
rect 1341 2677 1363 2683
rect 1357 2544 1363 2677
rect 1373 2664 1379 2676
rect 1437 2664 1443 2876
rect 1453 2804 1459 3296
rect 1485 3203 1491 3357
rect 1501 3304 1507 3316
rect 1517 3304 1523 3316
rect 1517 3204 1523 3296
rect 1485 3197 1507 3203
rect 1469 3064 1475 3196
rect 1501 3183 1507 3197
rect 1501 3177 1523 3183
rect 1485 3144 1491 3176
rect 1517 3124 1523 3177
rect 1533 3144 1539 3336
rect 1549 3264 1555 3436
rect 1565 3404 1571 3476
rect 1565 3243 1571 3356
rect 1581 3324 1587 3496
rect 1613 3484 1619 3576
rect 1597 3364 1603 3476
rect 1629 3463 1635 3556
rect 1661 3484 1667 3496
rect 1613 3457 1635 3463
rect 1613 3344 1619 3457
rect 1645 3423 1651 3476
rect 1645 3417 1667 3423
rect 1549 3237 1571 3243
rect 1549 3163 1555 3237
rect 1576 3206 1577 3214
rect 1585 3206 1587 3214
rect 1595 3206 1597 3214
rect 1605 3206 1607 3214
rect 1615 3206 1624 3214
rect 1645 3183 1651 3396
rect 1661 3344 1667 3417
rect 1661 3264 1667 3316
rect 1677 3304 1683 3716
rect 1709 3703 1715 3757
rect 1725 3724 1731 3736
rect 1693 3697 1715 3703
rect 1693 3584 1699 3697
rect 1741 3684 1747 3776
rect 1805 3744 1811 3857
rect 1885 3843 1891 3916
rect 1901 3884 1907 3957
rect 1885 3837 1907 3843
rect 1885 3763 1891 3796
rect 1901 3784 1907 3837
rect 1917 3804 1923 4176
rect 2029 4164 2035 4177
rect 1933 4124 1939 4136
rect 1949 4044 1955 4096
rect 1965 3924 1971 4116
rect 1981 3863 1987 4016
rect 2013 3924 2019 4036
rect 2029 3924 2035 3976
rect 2061 3924 2067 4516
rect 2077 4004 2083 4576
rect 2093 4304 2099 4376
rect 2125 4304 2131 4316
rect 2157 4223 2163 4643
rect 2237 4637 2259 4643
rect 2173 4344 2179 4536
rect 2173 4324 2179 4336
rect 2141 4217 2163 4223
rect 2141 4083 2147 4217
rect 2173 4164 2179 4316
rect 2205 4284 2211 4336
rect 2253 4283 2259 4637
rect 2461 4624 2467 4643
rect 2429 4577 2444 4583
rect 2397 4544 2403 4576
rect 2429 4564 2435 4577
rect 2445 4544 2451 4576
rect 2301 4504 2307 4516
rect 2317 4504 2323 4516
rect 2237 4277 2259 4283
rect 2157 4104 2163 4116
rect 2141 4077 2163 4083
rect 1997 3884 2003 3896
rect 2093 3884 2099 4016
rect 2052 3877 2067 3883
rect 2061 3864 2067 3877
rect 1981 3857 2003 3863
rect 1981 3804 1987 3836
rect 1885 3757 1907 3763
rect 1828 3737 1852 3743
rect 1693 3504 1699 3536
rect 1709 3423 1715 3676
rect 1805 3623 1811 3716
rect 1805 3617 1827 3623
rect 1773 3523 1779 3536
rect 1757 3517 1779 3523
rect 1757 3484 1763 3517
rect 1725 3464 1731 3476
rect 1789 3444 1795 3476
rect 1709 3417 1731 3423
rect 1709 3364 1715 3396
rect 1725 3363 1731 3417
rect 1805 3363 1811 3456
rect 1821 3404 1827 3617
rect 1837 3584 1843 3716
rect 1853 3584 1859 3696
rect 1869 3523 1875 3696
rect 1885 3684 1891 3716
rect 1901 3624 1907 3757
rect 1917 3704 1923 3756
rect 1997 3744 2003 3857
rect 2109 3844 2115 3876
rect 2125 3823 2131 4036
rect 2157 3984 2163 4077
rect 2221 3963 2227 4076
rect 2237 3984 2243 4277
rect 2253 3984 2259 4196
rect 2221 3957 2243 3963
rect 2205 3904 2211 3956
rect 2109 3817 2131 3823
rect 2029 3764 2035 3816
rect 1892 3557 1923 3563
rect 1917 3544 1923 3557
rect 1837 3517 1875 3523
rect 1837 3484 1843 3517
rect 1869 3463 1875 3517
rect 1853 3457 1875 3463
rect 1837 3444 1843 3456
rect 1821 3384 1827 3396
rect 1725 3357 1747 3363
rect 1805 3357 1827 3363
rect 1709 3337 1724 3343
rect 1629 3177 1651 3183
rect 1549 3157 1580 3163
rect 1549 3124 1555 3157
rect 1501 3083 1507 3116
rect 1517 3104 1523 3116
rect 1540 3097 1555 3103
rect 1549 3084 1555 3097
rect 1501 3077 1516 3083
rect 1533 3064 1539 3076
rect 1501 2984 1507 3056
rect 1485 2923 1491 2936
rect 1485 2917 1507 2923
rect 1501 2904 1507 2917
rect 1453 2704 1459 2776
rect 1373 2524 1379 2636
rect 1389 2544 1395 2576
rect 1405 2544 1411 2636
rect 1421 2523 1427 2636
rect 1421 2517 1436 2523
rect 1165 2377 1187 2383
rect 1165 2284 1171 2377
rect 1277 2363 1283 2516
rect 1309 2464 1315 2516
rect 1389 2484 1395 2516
rect 1405 2463 1411 2476
rect 1421 2464 1427 2476
rect 1389 2457 1411 2463
rect 1373 2384 1379 2456
rect 1389 2383 1395 2457
rect 1405 2404 1411 2436
rect 1421 2384 1427 2396
rect 1389 2377 1411 2383
rect 1229 2357 1283 2363
rect 1165 2124 1171 2276
rect 1197 2184 1203 2336
rect 1213 2204 1219 2296
rect 1229 2143 1235 2357
rect 1405 2363 1411 2377
rect 1316 2357 1363 2363
rect 1405 2357 1427 2363
rect 1357 2343 1363 2357
rect 1252 2337 1347 2343
rect 1357 2337 1411 2343
rect 1245 2264 1251 2336
rect 1341 2324 1347 2337
rect 1405 2324 1411 2337
rect 1277 2284 1283 2316
rect 1325 2304 1331 2316
rect 1389 2304 1395 2316
rect 1421 2303 1427 2357
rect 1405 2297 1427 2303
rect 1261 2184 1267 2196
rect 1261 2164 1267 2176
rect 1229 2137 1244 2143
rect 1325 2143 1331 2176
rect 1357 2144 1363 2276
rect 1389 2144 1395 2276
rect 1405 2184 1411 2297
rect 1421 2163 1427 2276
rect 1437 2264 1443 2496
rect 1453 2484 1459 2696
rect 1485 2684 1491 2896
rect 1501 2664 1507 2836
rect 1517 2804 1523 3036
rect 1565 2943 1571 3076
rect 1581 3024 1587 3136
rect 1549 2937 1571 2943
rect 1597 2943 1603 3096
rect 1613 3064 1619 3156
rect 1629 3084 1635 3177
rect 1645 3064 1651 3096
rect 1661 3084 1667 3196
rect 1693 3184 1699 3216
rect 1709 3184 1715 3337
rect 1741 3324 1747 3357
rect 1821 3324 1827 3357
rect 1709 3124 1715 3176
rect 1693 3064 1699 3116
rect 1629 3057 1644 3063
rect 1613 2964 1619 3036
rect 1597 2937 1619 2943
rect 1533 2783 1539 2896
rect 1549 2824 1555 2937
rect 1565 2863 1571 2896
rect 1597 2863 1603 2916
rect 1613 2864 1619 2937
rect 1629 2924 1635 3057
rect 1709 3044 1715 3116
rect 1725 3084 1731 3216
rect 1741 3104 1747 3316
rect 1789 3144 1795 3216
rect 1821 3144 1827 3256
rect 1837 3184 1843 3396
rect 1853 3364 1859 3457
rect 1869 3144 1875 3396
rect 1885 3383 1891 3536
rect 1933 3524 1939 3736
rect 2013 3704 2019 3736
rect 1949 3524 1955 3556
rect 1965 3523 1971 3696
rect 1965 3517 1987 3523
rect 1901 3444 1907 3476
rect 1917 3423 1923 3516
rect 1901 3417 1923 3423
rect 1933 3497 1964 3503
rect 1901 3404 1907 3417
rect 1885 3377 1900 3383
rect 1933 3364 1939 3497
rect 1949 3443 1955 3476
rect 1949 3437 1971 3443
rect 1965 3343 1971 3437
rect 1981 3364 1987 3517
rect 1892 3337 1907 3343
rect 1901 3264 1907 3337
rect 1933 3337 1971 3343
rect 1933 3264 1939 3337
rect 1972 3317 1987 3323
rect 1901 3184 1907 3256
rect 1901 3124 1907 3136
rect 1748 3077 1756 3083
rect 1661 2944 1667 3036
rect 1741 2983 1747 3056
rect 1725 2977 1747 2983
rect 1725 2964 1731 2977
rect 1668 2937 1683 2943
rect 1629 2903 1635 2916
rect 1629 2897 1651 2903
rect 1565 2857 1603 2863
rect 1576 2806 1577 2814
rect 1585 2806 1587 2814
rect 1595 2806 1597 2814
rect 1605 2806 1607 2814
rect 1615 2806 1624 2814
rect 1533 2777 1555 2783
rect 1549 2763 1555 2777
rect 1549 2757 1571 2763
rect 1517 2724 1523 2736
rect 1453 2424 1459 2456
rect 1453 2244 1459 2316
rect 1421 2157 1443 2163
rect 1325 2137 1347 2143
rect 1181 2124 1187 2136
rect 1341 2124 1347 2137
rect 1092 2117 1107 2123
rect 973 1924 979 1956
rect 685 1724 691 1736
rect 685 1704 691 1716
rect 733 1684 739 1716
rect 628 1537 643 1543
rect 541 1483 547 1516
rect 525 1477 547 1483
rect 413 1464 419 1476
rect 413 1364 419 1456
rect 381 1357 396 1363
rect 301 1184 307 1236
rect 285 1164 291 1176
rect 13 1104 19 1116
rect 221 1104 227 1116
rect 77 1064 83 1076
rect 125 1064 131 1096
rect 173 1064 179 1096
rect 317 1064 323 1096
rect 381 1084 387 1357
rect 445 1324 451 1356
rect 413 1164 419 1316
rect 45 984 51 1056
rect 93 1024 99 1036
rect 77 984 83 1016
rect 125 984 131 1056
rect 173 1044 179 1056
rect 317 1044 323 1056
rect 173 984 179 1036
rect 333 1004 339 1036
rect 349 984 355 1036
rect 381 943 387 1056
rect 397 944 403 956
rect 365 937 387 943
rect 61 904 67 936
rect 93 904 99 936
rect 205 904 211 916
rect 45 704 51 876
rect 93 704 99 896
rect 157 784 163 896
rect 189 784 195 876
rect 237 784 243 896
rect 253 784 259 856
rect 45 684 51 696
rect 45 383 51 676
rect 125 664 131 676
rect 221 664 227 676
rect 301 664 307 936
rect 317 824 323 916
rect 333 784 339 796
rect 349 704 355 816
rect 365 804 371 937
rect 413 924 419 1156
rect 493 1144 499 1436
rect 525 1363 531 1477
rect 580 1477 595 1483
rect 573 1384 579 1436
rect 509 1357 531 1363
rect 509 1344 515 1357
rect 589 1344 595 1477
rect 605 1444 611 1496
rect 637 1463 643 1537
rect 637 1457 652 1463
rect 605 1404 611 1436
rect 621 1344 627 1436
rect 637 1384 643 1457
rect 653 1344 659 1356
rect 685 1344 691 1496
rect 717 1483 723 1656
rect 765 1584 771 1716
rect 781 1684 787 1756
rect 749 1524 755 1576
rect 781 1564 787 1676
rect 797 1664 803 1756
rect 813 1724 819 1736
rect 733 1504 739 1516
rect 797 1484 803 1496
rect 701 1477 723 1483
rect 701 1444 707 1477
rect 733 1463 739 1476
rect 733 1457 755 1463
rect 749 1364 755 1457
rect 765 1364 771 1416
rect 557 1297 572 1303
rect 557 1224 563 1297
rect 589 1223 595 1336
rect 589 1217 611 1223
rect 493 1104 499 1136
rect 429 1064 435 1076
rect 397 897 451 903
rect 397 884 403 897
rect 429 824 435 836
rect 445 724 451 897
rect 349 684 355 696
rect 445 684 451 696
rect 413 664 419 676
rect 109 624 115 636
rect 141 504 147 536
rect 77 444 83 500
rect 36 377 51 383
rect 285 320 291 376
rect 77 108 83 296
rect 189 203 195 256
rect 173 197 195 203
rect 173 164 179 197
rect 77 97 83 100
rect 141 24 147 136
rect 301 124 307 656
rect 349 644 355 656
rect 349 564 355 636
rect 365 564 371 636
rect 381 584 387 596
rect 413 584 419 656
rect 429 644 435 656
rect 461 624 467 1076
rect 493 964 499 1056
rect 477 924 483 936
rect 477 644 483 896
rect 493 824 499 916
rect 509 864 515 1136
rect 525 1104 531 1116
rect 557 1064 563 1136
rect 589 1124 595 1136
rect 605 1104 611 1217
rect 589 1083 595 1096
rect 589 1077 604 1083
rect 573 1024 579 1076
rect 605 1024 611 1076
rect 637 1064 643 1116
rect 621 1004 627 1056
rect 621 963 627 996
rect 605 957 627 963
rect 525 944 531 956
rect 525 897 540 903
rect 509 784 515 816
rect 525 724 531 897
rect 557 884 563 956
rect 605 903 611 957
rect 637 943 643 1036
rect 653 943 659 1316
rect 669 1144 675 1156
rect 685 1144 691 1156
rect 701 1144 707 1256
rect 717 1244 723 1356
rect 749 1344 755 1356
rect 733 1204 739 1236
rect 669 1064 675 1136
rect 701 1124 707 1136
rect 637 937 659 943
rect 653 924 659 937
rect 605 897 620 903
rect 685 884 691 1096
rect 717 1064 723 1176
rect 765 1163 771 1296
rect 740 1157 771 1163
rect 733 1144 739 1156
rect 733 984 739 1116
rect 749 1104 755 1136
rect 765 1124 771 1136
rect 781 1124 787 1416
rect 813 1344 819 1556
rect 829 1484 835 1656
rect 845 1464 851 1496
rect 829 1424 835 1456
rect 861 1444 867 1716
rect 877 1624 883 1716
rect 893 1664 899 1896
rect 957 1624 963 1836
rect 989 1784 995 2056
rect 1021 1963 1027 2036
rect 1005 1957 1027 1963
rect 1005 1884 1011 1957
rect 1021 1904 1027 1936
rect 1037 1784 1043 2076
rect 1069 2004 1075 2116
rect 1101 2084 1107 2117
rect 1373 2117 1388 2123
rect 1197 2084 1203 2096
rect 1085 1983 1091 1996
rect 1149 1984 1155 1996
rect 1053 1977 1091 1983
rect 1053 1864 1059 1977
rect 1069 1864 1075 1876
rect 1053 1763 1059 1856
rect 1085 1824 1091 1956
rect 1165 1944 1171 2076
rect 1213 2024 1219 2076
rect 1229 2003 1235 2116
rect 1325 2083 1331 2116
rect 1373 2084 1379 2117
rect 1309 2077 1331 2083
rect 1213 1997 1235 2003
rect 1101 1937 1155 1943
rect 1101 1904 1107 1937
rect 1133 1904 1139 1916
rect 1149 1903 1155 1937
rect 1149 1897 1171 1903
rect 1101 1784 1107 1856
rect 1133 1824 1139 1876
rect 1053 1757 1075 1763
rect 1037 1704 1043 1716
rect 1037 1564 1043 1656
rect 1053 1583 1059 1636
rect 1069 1624 1075 1757
rect 1149 1624 1155 1876
rect 1165 1744 1171 1897
rect 1197 1804 1203 1836
rect 1213 1804 1219 1997
rect 1245 1964 1251 1996
rect 1277 1964 1283 1996
rect 1229 1937 1276 1943
rect 1229 1904 1235 1937
rect 1309 1943 1315 2077
rect 1405 2024 1411 2156
rect 1437 2143 1443 2157
rect 1437 2137 1459 2143
rect 1453 2104 1459 2137
rect 1469 2063 1475 2636
rect 1501 2484 1507 2636
rect 1517 2504 1523 2576
rect 1533 2524 1539 2756
rect 1565 2744 1571 2757
rect 1645 2744 1651 2897
rect 1677 2864 1683 2937
rect 1549 2704 1555 2736
rect 1549 2544 1555 2676
rect 1565 2584 1571 2696
rect 1597 2664 1603 2716
rect 1629 2697 1644 2703
rect 1613 2644 1619 2696
rect 1597 2564 1603 2636
rect 1485 2404 1491 2476
rect 1517 2444 1523 2476
rect 1501 2364 1507 2436
rect 1533 2384 1539 2476
rect 1517 2344 1523 2376
rect 1485 2324 1491 2336
rect 1501 2263 1507 2296
rect 1549 2284 1555 2536
rect 1629 2484 1635 2697
rect 1661 2684 1667 2856
rect 1677 2764 1683 2816
rect 1693 2804 1699 2936
rect 1757 2904 1763 3016
rect 1773 2964 1779 3076
rect 1789 3064 1795 3116
rect 1805 3043 1811 3116
rect 1853 3064 1859 3076
rect 1869 3064 1875 3116
rect 1885 3084 1891 3116
rect 1789 3037 1811 3043
rect 1789 2944 1795 3037
rect 1709 2843 1715 2856
rect 1709 2837 1731 2843
rect 1677 2704 1683 2716
rect 1693 2664 1699 2676
rect 1725 2644 1731 2837
rect 1757 2724 1763 2776
rect 1773 2744 1779 2876
rect 1789 2824 1795 2916
rect 1805 2824 1811 2936
rect 1821 2924 1827 3036
rect 1837 2984 1843 3036
rect 1869 2983 1875 2996
rect 1853 2977 1875 2983
rect 1853 2963 1859 2977
rect 1837 2957 1859 2963
rect 1837 2864 1843 2957
rect 1860 2937 1875 2943
rect 1869 2924 1875 2937
rect 1885 2884 1891 3076
rect 1917 3063 1923 3236
rect 1933 3184 1939 3216
rect 1965 3144 1971 3256
rect 1933 3104 1939 3136
rect 1981 3124 1987 3317
rect 1997 3144 2003 3536
rect 2013 3524 2019 3616
rect 2029 3544 2035 3716
rect 2029 3323 2035 3456
rect 2045 3364 2051 3516
rect 2061 3504 2067 3616
rect 2077 3524 2083 3776
rect 2109 3724 2115 3817
rect 2109 3664 2115 3696
rect 2093 3564 2099 3636
rect 2109 3584 2115 3596
rect 2125 3524 2131 3736
rect 2141 3503 2147 3876
rect 2189 3864 2195 3896
rect 2157 3744 2163 3856
rect 2157 3584 2163 3716
rect 2157 3504 2163 3556
rect 2125 3497 2147 3503
rect 2077 3484 2083 3496
rect 2109 3464 2115 3476
rect 2125 3443 2131 3497
rect 2173 3503 2179 3656
rect 2189 3584 2195 3776
rect 2205 3504 2211 3576
rect 2173 3497 2195 3503
rect 2109 3437 2131 3443
rect 2061 3324 2067 3436
rect 2109 3423 2115 3437
rect 2077 3417 2115 3423
rect 2077 3404 2083 3417
rect 2125 3403 2131 3416
rect 2125 3397 2179 3403
rect 2173 3384 2179 3397
rect 2189 3363 2195 3497
rect 2173 3357 2195 3363
rect 2013 3317 2035 3323
rect 2013 3204 2019 3317
rect 2093 3323 2099 3356
rect 2109 3344 2115 3356
rect 2173 3343 2179 3357
rect 2164 3337 2179 3343
rect 2093 3317 2115 3323
rect 2036 3297 2044 3303
rect 2068 3297 2092 3303
rect 2109 3303 2115 3317
rect 2109 3297 2131 3303
rect 1933 3084 1939 3096
rect 2029 3084 2035 3136
rect 2061 3124 2067 3256
rect 1917 3057 1939 3063
rect 1901 2924 1907 2996
rect 1933 2964 1939 3057
rect 1965 2963 1971 3056
rect 1981 3043 1987 3076
rect 2029 3057 2044 3063
rect 2029 3044 2035 3057
rect 1981 3037 2003 3043
rect 1997 3024 2003 3037
rect 1981 2984 1987 3016
rect 2045 3004 2051 3036
rect 1965 2957 1987 2963
rect 1853 2823 1859 2876
rect 1837 2817 1859 2823
rect 1789 2783 1795 2816
rect 1805 2804 1811 2816
rect 1789 2777 1811 2783
rect 1805 2764 1811 2777
rect 1789 2704 1795 2756
rect 1757 2697 1772 2703
rect 1661 2424 1667 2556
rect 1693 2544 1699 2556
rect 1757 2544 1763 2697
rect 1773 2544 1779 2676
rect 1805 2664 1811 2676
rect 1821 2644 1827 2716
rect 1677 2524 1683 2536
rect 1576 2406 1577 2414
rect 1585 2406 1587 2414
rect 1595 2406 1597 2414
rect 1605 2406 1607 2414
rect 1615 2406 1624 2414
rect 1581 2284 1587 2356
rect 1501 2257 1523 2263
rect 1517 2223 1523 2257
rect 1581 2223 1587 2236
rect 1517 2217 1587 2223
rect 1549 2157 1587 2163
rect 1501 2124 1507 2156
rect 1549 2123 1555 2157
rect 1581 2144 1587 2157
rect 1645 2144 1651 2396
rect 1693 2304 1699 2516
rect 1725 2503 1731 2536
rect 1709 2497 1731 2503
rect 1709 2424 1715 2497
rect 1693 2284 1699 2296
rect 1709 2284 1715 2316
rect 1757 2303 1763 2436
rect 1741 2297 1763 2303
rect 1677 2264 1683 2276
rect 1661 2243 1667 2256
rect 1741 2243 1747 2297
rect 1661 2237 1747 2243
rect 1716 2157 1724 2163
rect 1741 2143 1747 2156
rect 1741 2137 1763 2143
rect 1517 2117 1555 2123
rect 1517 2104 1523 2117
rect 1533 2097 1571 2103
rect 1533 2084 1539 2097
rect 1565 2083 1571 2097
rect 1597 2083 1603 2096
rect 1565 2077 1603 2083
rect 1469 2057 1491 2063
rect 1469 2024 1475 2036
rect 1341 2004 1347 2016
rect 1485 2004 1491 2057
rect 1576 2006 1577 2014
rect 1585 2006 1587 2014
rect 1595 2006 1597 2014
rect 1605 2006 1607 2014
rect 1615 2006 1624 2014
rect 1341 1963 1347 1996
rect 1357 1984 1363 1996
rect 1332 1957 1347 1963
rect 1309 1937 1331 1943
rect 1245 1884 1251 1916
rect 1325 1904 1331 1937
rect 1373 1904 1379 1996
rect 1517 1924 1523 1996
rect 1645 1944 1651 2096
rect 1661 2024 1667 2096
rect 1661 1984 1667 1996
rect 1693 1984 1699 2056
rect 1245 1824 1251 1876
rect 1261 1844 1267 1876
rect 1277 1823 1283 1896
rect 1309 1863 1315 1876
rect 1309 1857 1331 1863
rect 1261 1817 1283 1823
rect 1188 1717 1203 1723
rect 1053 1577 1091 1583
rect 1085 1543 1091 1577
rect 1197 1563 1203 1717
rect 1181 1557 1203 1563
rect 1085 1537 1107 1543
rect 989 1524 995 1536
rect 877 1504 883 1516
rect 1021 1504 1027 1536
rect 1085 1504 1091 1516
rect 1101 1504 1107 1537
rect 877 1443 883 1476
rect 877 1437 899 1443
rect 765 1097 780 1103
rect 765 1043 771 1097
rect 765 1037 787 1043
rect 749 904 755 936
rect 605 823 611 876
rect 589 817 611 823
rect 589 684 595 817
rect 621 724 627 876
rect 669 864 675 876
rect 637 724 643 856
rect 669 724 675 856
rect 685 724 691 876
rect 717 784 723 836
rect 749 824 755 836
rect 749 803 755 816
rect 765 804 771 936
rect 781 824 787 1037
rect 797 984 803 1316
rect 813 1224 819 1296
rect 829 1104 835 1236
rect 845 1084 851 1136
rect 845 1064 851 1076
rect 861 1004 867 1416
rect 877 1324 883 1416
rect 893 1324 899 1437
rect 957 1384 963 1476
rect 989 1464 995 1496
rect 941 1344 947 1376
rect 973 1344 979 1376
rect 989 1324 995 1436
rect 1037 1424 1043 1496
rect 1021 1364 1027 1416
rect 1053 1404 1059 1496
rect 1069 1344 1075 1476
rect 1133 1423 1139 1476
rect 1133 1417 1155 1423
rect 1021 1323 1027 1336
rect 1085 1324 1091 1336
rect 1021 1317 1043 1323
rect 893 1203 899 1296
rect 925 1204 931 1296
rect 1037 1283 1043 1317
rect 1037 1277 1059 1283
rect 1053 1264 1059 1277
rect 989 1237 1059 1243
rect 893 1197 915 1203
rect 909 1124 915 1197
rect 948 1117 956 1123
rect 973 1103 979 1196
rect 989 1144 995 1237
rect 957 1097 979 1103
rect 836 997 851 1003
rect 829 904 835 916
rect 733 797 755 803
rect 717 684 723 736
rect 733 704 739 797
rect 797 723 803 896
rect 813 824 819 896
rect 813 784 819 816
rect 845 784 851 997
rect 861 944 867 956
rect 877 944 883 1056
rect 893 943 899 996
rect 909 984 915 1096
rect 941 1044 947 1076
rect 957 1004 963 1097
rect 989 1084 995 1116
rect 989 1024 995 1076
rect 1005 1003 1011 1216
rect 1037 1124 1043 1216
rect 1053 1144 1059 1237
rect 1069 1184 1075 1296
rect 1085 1163 1091 1296
rect 1101 1244 1107 1336
rect 1117 1304 1123 1416
rect 1133 1384 1139 1396
rect 1149 1344 1155 1417
rect 1165 1344 1171 1516
rect 1181 1483 1187 1557
rect 1229 1544 1235 1816
rect 1261 1803 1267 1817
rect 1245 1797 1267 1803
rect 1245 1744 1251 1797
rect 1245 1624 1251 1716
rect 1197 1524 1203 1536
rect 1245 1524 1251 1596
rect 1261 1524 1267 1636
rect 1277 1624 1283 1796
rect 1293 1784 1299 1856
rect 1325 1843 1331 1857
rect 1325 1837 1379 1843
rect 1325 1704 1331 1716
rect 1341 1704 1347 1816
rect 1357 1783 1363 1816
rect 1373 1804 1379 1837
rect 1389 1824 1395 1876
rect 1405 1803 1411 1856
rect 1437 1843 1443 1876
rect 1453 1863 1459 1896
rect 1613 1884 1619 1916
rect 1677 1904 1683 1956
rect 1709 1924 1715 2136
rect 1725 1924 1731 2136
rect 1741 2083 1747 2116
rect 1757 2104 1763 2137
rect 1773 2083 1779 2516
rect 1789 2364 1795 2516
rect 1789 2264 1795 2296
rect 1805 2184 1811 2636
rect 1837 2624 1843 2817
rect 1917 2724 1923 2956
rect 1933 2704 1939 2876
rect 1949 2824 1955 2936
rect 1853 2684 1859 2696
rect 1821 2544 1827 2616
rect 1853 2603 1859 2676
rect 1885 2644 1891 2696
rect 1917 2684 1923 2696
rect 1949 2684 1955 2816
rect 1901 2664 1907 2676
rect 1837 2597 1859 2603
rect 1821 2463 1827 2516
rect 1837 2504 1843 2597
rect 1901 2564 1907 2656
rect 1853 2484 1859 2556
rect 1869 2544 1875 2556
rect 1885 2524 1891 2536
rect 1821 2457 1875 2463
rect 1821 2384 1827 2436
rect 1869 2364 1875 2457
rect 1885 2384 1891 2436
rect 1933 2424 1939 2536
rect 1949 2504 1955 2616
rect 1853 2304 1859 2356
rect 1933 2324 1939 2336
rect 1885 2283 1891 2316
rect 1949 2303 1955 2376
rect 1965 2344 1971 2576
rect 1981 2544 1987 2957
rect 1997 2884 2003 2936
rect 1997 2844 2003 2876
rect 1997 2704 2003 2796
rect 2013 2784 2019 2836
rect 1997 2564 2003 2676
rect 2013 2584 2019 2696
rect 2029 2624 2035 2956
rect 2045 2844 2051 2896
rect 2061 2823 2067 3096
rect 2077 3064 2083 3116
rect 2093 3104 2099 3236
rect 2077 3004 2083 3036
rect 2045 2817 2067 2823
rect 2045 2724 2051 2817
rect 2077 2803 2083 2916
rect 2093 2904 2099 3056
rect 2109 2944 2115 3276
rect 2125 3124 2131 3297
rect 2141 3224 2147 3256
rect 2157 3164 2163 3296
rect 2173 3064 2179 3337
rect 2189 3324 2195 3336
rect 2205 3224 2211 3316
rect 2221 3304 2227 3816
rect 2237 3604 2243 3957
rect 2253 3864 2259 3916
rect 2269 3703 2275 4436
rect 2301 4424 2307 4496
rect 2397 4444 2403 4536
rect 2301 4324 2307 4416
rect 2333 4384 2339 4436
rect 2413 4403 2419 4436
rect 2397 4397 2419 4403
rect 2285 4304 2291 4316
rect 2285 4184 2291 4296
rect 2301 4284 2307 4296
rect 2397 4284 2403 4397
rect 2317 4264 2323 4276
rect 2397 4237 2412 4243
rect 2381 4204 2387 4236
rect 2397 4104 2403 4237
rect 2413 4124 2419 4216
rect 2429 4164 2435 4276
rect 2317 3957 2387 3963
rect 2317 3943 2323 3957
rect 2381 3944 2387 3957
rect 2285 3937 2323 3943
rect 2285 3884 2291 3937
rect 2340 3937 2364 3943
rect 2413 3943 2419 4116
rect 2461 4083 2467 4376
rect 2493 4164 2499 4176
rect 2509 4143 2515 4643
rect 2637 4584 2643 4643
rect 2749 4624 2755 4643
rect 2797 4584 2803 4643
rect 2861 4584 2867 4643
rect 2909 4624 2915 4643
rect 3069 4637 3123 4643
rect 3069 4584 3075 4637
rect 3245 4624 3251 4643
rect 3309 4624 3315 4643
rect 3501 4624 3507 4643
rect 3028 4577 3043 4583
rect 3037 4564 3043 4577
rect 2557 4344 2563 4536
rect 2573 4526 2579 4556
rect 2573 4517 2579 4518
rect 2772 4517 2780 4523
rect 2717 4504 2723 4516
rect 2813 4384 2819 4516
rect 2893 4384 2899 4496
rect 2557 4304 2563 4336
rect 2525 4244 2531 4296
rect 2637 4264 2643 4336
rect 2685 4304 2691 4356
rect 2733 4304 2739 4376
rect 2909 4344 2915 4536
rect 2925 4324 2931 4556
rect 2957 4384 2963 4536
rect 2829 4304 2835 4316
rect 2500 4137 2515 4143
rect 2564 4137 2627 4143
rect 2493 4117 2547 4123
rect 2493 4104 2499 4117
rect 2541 4104 2547 4117
rect 2621 4123 2627 4137
rect 2621 4117 2668 4123
rect 2557 4104 2563 4116
rect 2605 4104 2611 4116
rect 2701 4104 2707 4256
rect 2461 4077 2483 4083
rect 2397 3937 2419 3943
rect 2397 3924 2403 3937
rect 2317 3864 2323 3896
rect 2253 3697 2275 3703
rect 2253 3463 2259 3697
rect 2285 3464 2291 3836
rect 2333 3664 2339 3916
rect 2429 3904 2435 3936
rect 2388 3897 2396 3903
rect 2397 3844 2403 3876
rect 2349 3784 2355 3836
rect 2365 3804 2371 3836
rect 2413 3784 2419 3856
rect 2429 3784 2435 3876
rect 2445 3864 2451 4016
rect 2477 3963 2483 4077
rect 2500 4077 2515 4083
rect 2509 3984 2515 4077
rect 2525 3984 2531 4096
rect 2557 4004 2563 4036
rect 2461 3957 2483 3963
rect 2461 3744 2467 3957
rect 2493 3924 2499 3956
rect 2477 3884 2483 3896
rect 2541 3744 2547 3996
rect 2605 3904 2611 4036
rect 2557 3864 2563 3876
rect 2237 3457 2259 3463
rect 2237 3103 2243 3457
rect 2301 3424 2307 3616
rect 2333 3504 2339 3536
rect 2269 3343 2275 3416
rect 2253 3337 2275 3343
rect 2253 3324 2259 3337
rect 2301 3324 2307 3396
rect 2317 3343 2323 3456
rect 2333 3384 2339 3456
rect 2349 3404 2355 3736
rect 2429 3684 2435 3696
rect 2381 3524 2387 3576
rect 2397 3557 2428 3563
rect 2397 3544 2403 3557
rect 2445 3544 2451 3716
rect 2461 3704 2467 3716
rect 2429 3504 2435 3536
rect 2461 3524 2467 3596
rect 2381 3384 2387 3396
rect 2349 3344 2355 3376
rect 2365 3364 2371 3376
rect 2365 3344 2371 3356
rect 2317 3337 2339 3343
rect 2269 3303 2275 3316
rect 2260 3297 2275 3303
rect 2317 3283 2323 3316
rect 2333 3304 2339 3337
rect 2317 3277 2355 3283
rect 2349 3263 2355 3277
rect 2349 3257 2364 3263
rect 2285 3164 2291 3256
rect 2333 3184 2339 3256
rect 2397 3184 2403 3356
rect 2429 3344 2435 3476
rect 2285 3124 2291 3156
rect 2237 3097 2259 3103
rect 2141 3004 2147 3056
rect 2157 3003 2163 3036
rect 2189 3004 2195 3076
rect 2253 3064 2259 3097
rect 2269 3084 2275 3116
rect 2157 2997 2179 3003
rect 2109 2884 2115 2916
rect 2077 2797 2099 2803
rect 2093 2743 2099 2797
rect 2109 2763 2115 2836
rect 2125 2824 2131 2916
rect 2173 2904 2179 2997
rect 2205 2983 2211 2996
rect 2189 2977 2211 2983
rect 2189 2964 2195 2977
rect 2237 2964 2243 3016
rect 2253 2964 2259 3036
rect 2269 3024 2275 3036
rect 2157 2864 2163 2896
rect 2141 2784 2147 2856
rect 2157 2824 2163 2836
rect 2205 2824 2211 2956
rect 2109 2757 2131 2763
rect 2093 2737 2115 2743
rect 2109 2724 2115 2737
rect 2045 2664 2051 2716
rect 2125 2704 2131 2757
rect 2173 2703 2179 2716
rect 2157 2697 2179 2703
rect 2029 2597 2067 2603
rect 2029 2584 2035 2597
rect 2061 2584 2067 2597
rect 2045 2563 2051 2576
rect 2077 2563 2083 2696
rect 2093 2584 2099 2656
rect 2125 2624 2131 2676
rect 2141 2603 2147 2616
rect 2125 2597 2147 2603
rect 2029 2557 2051 2563
rect 2061 2557 2083 2563
rect 2013 2523 2019 2536
rect 1997 2517 2019 2523
rect 2029 2523 2035 2557
rect 2061 2544 2067 2557
rect 2029 2517 2044 2523
rect 1933 2297 1955 2303
rect 1885 2277 1923 2283
rect 1853 2244 1859 2256
rect 1837 2143 1843 2236
rect 1917 2224 1923 2277
rect 1933 2203 1939 2297
rect 1965 2244 1971 2256
rect 1917 2197 1939 2203
rect 1885 2144 1891 2196
rect 1821 2137 1843 2143
rect 1789 2104 1795 2116
rect 1741 2077 1763 2083
rect 1773 2077 1795 2083
rect 1757 2063 1763 2077
rect 1757 2057 1779 2063
rect 1757 1924 1763 1996
rect 1773 1984 1779 2057
rect 1652 1897 1667 1903
rect 1661 1883 1667 1897
rect 1709 1897 1724 1903
rect 1709 1883 1715 1897
rect 1661 1877 1715 1883
rect 1485 1863 1491 1876
rect 1549 1864 1555 1876
rect 1453 1857 1491 1863
rect 1437 1837 1459 1843
rect 1421 1804 1427 1836
rect 1389 1797 1411 1803
rect 1389 1783 1395 1797
rect 1437 1784 1443 1816
rect 1453 1804 1459 1837
rect 1501 1837 1516 1843
rect 1501 1823 1507 1837
rect 1533 1823 1539 1856
rect 1645 1844 1651 1876
rect 1661 1857 1692 1863
rect 1485 1817 1507 1823
rect 1517 1817 1539 1823
rect 1613 1817 1644 1823
rect 1357 1777 1395 1783
rect 1469 1763 1475 1816
rect 1485 1804 1491 1817
rect 1469 1757 1484 1763
rect 1389 1737 1484 1743
rect 1373 1724 1379 1736
rect 1373 1623 1379 1696
rect 1389 1643 1395 1737
rect 1389 1637 1411 1643
rect 1373 1617 1395 1623
rect 1293 1577 1308 1583
rect 1293 1563 1299 1577
rect 1325 1563 1331 1596
rect 1389 1584 1395 1617
rect 1277 1557 1299 1563
rect 1309 1557 1331 1563
rect 1277 1544 1283 1557
rect 1213 1484 1219 1496
rect 1229 1484 1235 1516
rect 1181 1477 1203 1483
rect 1149 1304 1155 1336
rect 1069 1157 1091 1163
rect 1021 1024 1027 1036
rect 989 997 1011 1003
rect 925 964 931 996
rect 893 937 908 943
rect 916 897 931 903
rect 925 763 931 897
rect 941 784 947 976
rect 973 963 979 996
rect 989 964 995 997
rect 1021 964 1027 976
rect 964 957 979 963
rect 989 944 995 956
rect 973 904 979 916
rect 989 883 995 896
rect 973 877 995 883
rect 957 763 963 876
rect 925 757 963 763
rect 797 717 812 723
rect 781 684 787 716
rect 861 703 867 736
rect 861 697 883 703
rect 525 644 531 656
rect 413 564 419 576
rect 445 564 451 616
rect 477 564 483 636
rect 509 624 515 636
rect 557 624 563 636
rect 573 544 579 676
rect 589 564 595 676
rect 605 484 611 656
rect 845 643 851 696
rect 845 637 867 643
rect 621 544 627 636
rect 621 484 627 516
rect 637 484 643 556
rect 669 544 675 636
rect 573 284 579 356
rect 333 184 339 196
rect 541 164 547 256
rect 653 224 659 536
rect 717 383 723 576
rect 733 424 739 556
rect 749 544 755 556
rect 813 544 819 556
rect 749 484 755 516
rect 765 484 771 516
rect 813 504 819 536
rect 717 377 732 383
rect 669 324 675 376
rect 781 144 787 496
rect 829 404 835 556
rect 845 504 851 616
rect 861 544 867 637
rect 861 524 867 536
rect 877 404 883 697
rect 909 564 915 756
rect 957 723 963 736
rect 941 717 963 723
rect 941 704 947 717
rect 973 664 979 877
rect 1037 804 1043 1076
rect 1069 964 1075 1157
rect 1085 1084 1091 1116
rect 1117 1064 1123 1216
rect 1133 1144 1139 1236
rect 1133 1084 1139 1116
rect 1149 1104 1155 1296
rect 1197 1264 1203 1477
rect 1229 1424 1235 1476
rect 1245 1304 1251 1496
rect 1293 1463 1299 1536
rect 1277 1457 1299 1463
rect 1261 1384 1267 1456
rect 1165 1084 1171 1096
rect 1101 1004 1107 1036
rect 1069 883 1075 936
rect 1053 877 1075 883
rect 1053 824 1059 877
rect 1069 803 1075 816
rect 1053 797 1075 803
rect 1053 724 1059 797
rect 1085 764 1091 956
rect 1117 944 1123 1036
rect 1133 1024 1139 1076
rect 1117 864 1123 896
rect 1021 717 1052 723
rect 989 704 995 716
rect 1005 683 1011 716
rect 1021 704 1027 717
rect 1085 684 1091 736
rect 1101 704 1107 796
rect 1133 784 1139 976
rect 1149 964 1155 1056
rect 1181 984 1187 1236
rect 1197 1104 1203 1116
rect 1213 1003 1219 1276
rect 1261 1204 1267 1336
rect 1277 1184 1283 1457
rect 1293 1384 1299 1436
rect 1309 1264 1315 1557
rect 1325 1324 1331 1536
rect 1405 1524 1411 1637
rect 1469 1524 1475 1596
rect 1485 1504 1491 1716
rect 1501 1524 1507 1796
rect 1517 1704 1523 1817
rect 1613 1764 1619 1817
rect 1661 1804 1667 1857
rect 1773 1844 1779 1876
rect 1789 1844 1795 2077
rect 1805 2004 1811 2136
rect 1821 2124 1827 2137
rect 1917 2123 1923 2197
rect 1901 2117 1923 2123
rect 1837 2024 1843 2036
rect 1805 1984 1811 1996
rect 1805 1864 1811 1896
rect 1629 1784 1635 1796
rect 1677 1764 1683 1836
rect 1693 1744 1699 1816
rect 1604 1717 1660 1723
rect 1549 1637 1564 1643
rect 1396 1497 1411 1503
rect 1341 1463 1347 1496
rect 1380 1477 1395 1483
rect 1389 1464 1395 1477
rect 1341 1457 1363 1463
rect 1245 1157 1315 1163
rect 1245 1144 1251 1157
rect 1309 1144 1315 1157
rect 1261 1124 1267 1136
rect 1325 1124 1331 1236
rect 1341 1143 1347 1436
rect 1357 1384 1363 1457
rect 1405 1424 1411 1497
rect 1357 1357 1372 1363
rect 1357 1264 1363 1357
rect 1421 1343 1427 1496
rect 1469 1423 1475 1496
rect 1517 1483 1523 1596
rect 1533 1524 1539 1616
rect 1549 1523 1555 1637
rect 1604 1637 1651 1643
rect 1645 1624 1651 1637
rect 1576 1606 1577 1614
rect 1585 1606 1587 1614
rect 1595 1606 1597 1614
rect 1605 1606 1607 1614
rect 1615 1606 1624 1614
rect 1645 1544 1651 1596
rect 1581 1537 1635 1543
rect 1549 1517 1571 1523
rect 1501 1477 1523 1483
rect 1437 1417 1475 1423
rect 1437 1364 1443 1417
rect 1485 1344 1491 1476
rect 1405 1337 1427 1343
rect 1373 1304 1379 1336
rect 1357 1184 1363 1236
rect 1341 1137 1363 1143
rect 1245 1104 1251 1116
rect 1261 1044 1267 1116
rect 1309 1104 1315 1116
rect 1197 997 1219 1003
rect 1197 963 1203 997
rect 1229 964 1235 1036
rect 1165 957 1203 963
rect 1165 944 1171 957
rect 1245 944 1251 976
rect 1165 883 1171 896
rect 1149 877 1171 883
rect 1149 764 1155 877
rect 1181 764 1187 856
rect 1197 804 1203 936
rect 1245 823 1251 936
rect 1277 924 1283 936
rect 1261 884 1267 896
rect 1229 817 1267 823
rect 1229 783 1235 817
rect 1197 777 1235 783
rect 1117 724 1123 736
rect 1165 684 1171 716
rect 1197 684 1203 777
rect 1245 724 1251 796
rect 1261 684 1267 817
rect 1277 744 1283 916
rect 1293 904 1299 1036
rect 1309 944 1315 1096
rect 1341 1084 1347 1116
rect 1341 1024 1347 1076
rect 1357 963 1363 1137
rect 1389 1104 1395 1336
rect 1405 1284 1411 1337
rect 1501 1304 1507 1477
rect 1517 1304 1523 1456
rect 1533 1344 1539 1456
rect 1549 1344 1555 1476
rect 1565 1464 1571 1517
rect 1565 1344 1571 1436
rect 1581 1384 1587 1537
rect 1597 1464 1603 1496
rect 1444 1297 1459 1303
rect 1437 1244 1443 1276
rect 1453 1244 1459 1297
rect 1469 1224 1475 1296
rect 1405 1104 1411 1196
rect 1373 984 1379 1016
rect 1421 1004 1427 1136
rect 1437 1104 1443 1136
rect 1485 1124 1491 1296
rect 1501 1144 1507 1296
rect 1517 1144 1523 1296
rect 1533 1284 1539 1316
rect 1549 1224 1555 1316
rect 1597 1304 1603 1416
rect 1613 1404 1619 1516
rect 1629 1404 1635 1537
rect 1661 1464 1667 1576
rect 1677 1524 1683 1736
rect 1709 1604 1715 1816
rect 1773 1743 1779 1836
rect 1837 1824 1843 1976
rect 1885 1964 1891 2116
rect 1901 2084 1907 2117
rect 1789 1763 1795 1816
rect 1821 1803 1827 1816
rect 1853 1803 1859 1816
rect 1821 1797 1859 1803
rect 1869 1784 1875 1956
rect 1917 1884 1923 2076
rect 1949 1904 1955 1976
rect 1965 1904 1971 2156
rect 1981 1984 1987 2276
rect 1997 2144 2003 2517
rect 2093 2504 2099 2556
rect 2125 2544 2131 2597
rect 2157 2583 2163 2697
rect 2189 2664 2195 2776
rect 2205 2723 2211 2816
rect 2221 2744 2227 2876
rect 2205 2717 2220 2723
rect 2205 2684 2211 2717
rect 2237 2683 2243 2936
rect 2269 2924 2275 2936
rect 2285 2844 2291 3056
rect 2301 3024 2307 3116
rect 2317 2964 2323 3156
rect 2381 3124 2387 3176
rect 2429 3164 2435 3316
rect 2445 3304 2451 3476
rect 2461 3303 2467 3496
rect 2477 3404 2483 3616
rect 2493 3484 2499 3676
rect 2509 3404 2515 3696
rect 2557 3604 2563 3716
rect 2573 3584 2579 3876
rect 2605 3864 2611 3896
rect 2621 3884 2627 4076
rect 2653 3984 2659 4076
rect 2669 3924 2675 3996
rect 2637 3863 2643 3916
rect 2637 3857 2659 3863
rect 2637 3804 2643 3836
rect 2525 3504 2531 3576
rect 2605 3564 2611 3796
rect 2541 3484 2547 3496
rect 2484 3337 2499 3343
rect 2493 3304 2499 3337
rect 2541 3323 2547 3376
rect 2557 3363 2563 3516
rect 2621 3504 2627 3536
rect 2637 3523 2643 3716
rect 2653 3544 2659 3857
rect 2669 3784 2675 3880
rect 2685 3864 2691 4096
rect 2717 4084 2723 4116
rect 2733 4103 2739 4296
rect 2781 4244 2787 4296
rect 2861 4224 2867 4296
rect 2813 4123 2819 4136
rect 2861 4124 2867 4136
rect 2877 4124 2883 4296
rect 2925 4244 2931 4296
rect 2909 4124 2915 4196
rect 2813 4117 2828 4123
rect 2733 4097 2764 4103
rect 2781 4084 2787 4116
rect 2893 4084 2899 4096
rect 2925 4084 2931 4196
rect 2941 4184 2947 4296
rect 2733 4043 2739 4076
rect 2717 4037 2739 4043
rect 2765 4037 2780 4043
rect 2717 3944 2723 4037
rect 2765 4023 2771 4037
rect 2797 4023 2803 4076
rect 2749 4017 2771 4023
rect 2781 4017 2803 4023
rect 2749 3984 2755 4017
rect 2669 3724 2675 3776
rect 2685 3744 2691 3776
rect 2701 3744 2707 3936
rect 2724 3917 2748 3923
rect 2749 3884 2755 3916
rect 2717 3864 2723 3876
rect 2733 3803 2739 3836
rect 2717 3797 2739 3803
rect 2685 3724 2691 3736
rect 2669 3684 2675 3696
rect 2637 3517 2659 3523
rect 2612 3477 2627 3483
rect 2573 3384 2579 3476
rect 2589 3384 2595 3476
rect 2605 3364 2611 3456
rect 2621 3384 2627 3477
rect 2557 3357 2595 3363
rect 2532 3317 2547 3323
rect 2461 3297 2476 3303
rect 2509 3303 2515 3316
rect 2557 3303 2563 3316
rect 2509 3297 2563 3303
rect 2445 3183 2451 3296
rect 2509 3277 2547 3283
rect 2509 3264 2515 3277
rect 2461 3224 2467 3236
rect 2493 3224 2499 3236
rect 2525 3183 2531 3256
rect 2445 3177 2467 3183
rect 2429 3124 2435 3136
rect 2413 3117 2428 3123
rect 2413 3104 2419 3117
rect 2397 3044 2403 3076
rect 2445 3044 2451 3156
rect 2461 3143 2467 3177
rect 2493 3177 2531 3183
rect 2541 3183 2547 3277
rect 2573 3203 2579 3336
rect 2589 3264 2595 3357
rect 2605 3304 2611 3336
rect 2605 3243 2611 3256
rect 2605 3237 2627 3243
rect 2573 3197 2604 3203
rect 2621 3183 2627 3237
rect 2653 3183 2659 3517
rect 2685 3504 2691 3716
rect 2701 3704 2707 3716
rect 2701 3623 2707 3676
rect 2717 3664 2723 3797
rect 2701 3617 2723 3623
rect 2717 3604 2723 3617
rect 2701 3584 2707 3596
rect 2733 3584 2739 3676
rect 2749 3464 2755 3756
rect 2765 3724 2771 3996
rect 2781 3944 2787 4017
rect 2781 3904 2787 3916
rect 2797 3903 2803 3956
rect 2813 3924 2819 4076
rect 2877 4063 2883 4076
rect 2909 4063 2915 4076
rect 2877 4057 2915 4063
rect 2861 3984 2867 4056
rect 2877 3984 2883 3996
rect 2877 3964 2883 3976
rect 2893 3904 2899 3996
rect 2797 3897 2819 3903
rect 2813 3884 2819 3897
rect 2909 3903 2915 4036
rect 2941 3904 2947 4116
rect 2957 4104 2963 4316
rect 2989 4264 2995 4296
rect 3021 4264 3027 4496
rect 2973 4163 2979 4256
rect 2989 4184 2995 4196
rect 2973 4157 2995 4163
rect 2973 4084 2979 4116
rect 2989 4083 2995 4157
rect 3037 4144 3043 4316
rect 3053 4264 3059 4456
rect 3053 4124 3059 4236
rect 3012 4117 3043 4123
rect 2989 4077 3011 4083
rect 2957 3944 2963 4076
rect 2973 4063 2979 4076
rect 2973 4057 2995 4063
rect 2909 3897 2931 3903
rect 2861 3884 2867 3896
rect 2925 3884 2931 3897
rect 2989 3884 2995 4057
rect 2781 3744 2787 3876
rect 2797 3784 2803 3876
rect 2909 3864 2915 3876
rect 2813 3744 2819 3756
rect 2861 3724 2867 3796
rect 2909 3764 2915 3856
rect 2925 3724 2931 3796
rect 2973 3724 2979 3836
rect 3005 3763 3011 4077
rect 3021 3884 3027 4096
rect 3037 4064 3043 4117
rect 3069 4104 3075 4556
rect 3085 4504 3091 4616
rect 3112 4606 3113 4614
rect 3121 4606 3123 4614
rect 3131 4606 3133 4614
rect 3141 4606 3143 4614
rect 3151 4606 3160 4614
rect 3517 4603 3523 4616
rect 3485 4597 3523 4603
rect 3357 4544 3363 4556
rect 3261 4524 3267 4536
rect 3101 4484 3107 4516
rect 3165 4484 3171 4516
rect 3117 4264 3123 4456
rect 3277 4344 3283 4536
rect 3364 4517 3372 4523
rect 3421 4504 3427 4516
rect 3112 4206 3113 4214
rect 3121 4206 3123 4214
rect 3131 4206 3133 4214
rect 3141 4206 3143 4214
rect 3151 4206 3160 4214
rect 3085 4104 3091 4116
rect 3101 4084 3107 4116
rect 3060 4077 3075 4083
rect 3069 4063 3075 4077
rect 3069 4057 3100 4063
rect 3117 3944 3123 4076
rect 3181 4044 3187 4316
rect 3277 4304 3283 4336
rect 3229 4284 3235 4296
rect 3213 4184 3219 4276
rect 3357 4264 3363 4336
rect 3373 4324 3379 4476
rect 3453 4464 3459 4536
rect 3485 4504 3491 4597
rect 3677 4577 3692 4583
rect 3677 4564 3683 4577
rect 4429 4577 4444 4583
rect 4093 4564 4099 4576
rect 4429 4564 4435 4577
rect 5933 4583 5939 4596
rect 6237 4584 6243 4596
rect 5917 4577 5939 4583
rect 4829 4564 4835 4576
rect 4813 4544 4819 4556
rect 3805 4504 3811 4516
rect 3533 4384 3539 4496
rect 3501 4304 3507 4316
rect 3549 4304 3555 4336
rect 3645 4324 3651 4416
rect 3229 4144 3235 4196
rect 3293 4184 3299 4216
rect 3229 4104 3235 4136
rect 2989 3757 3011 3763
rect 2781 3624 2787 3716
rect 2797 3697 2812 3703
rect 2797 3604 2803 3697
rect 2829 3624 2835 3656
rect 2877 3564 2883 3716
rect 2893 3684 2899 3696
rect 2973 3684 2979 3716
rect 2909 3624 2915 3676
rect 2909 3584 2915 3596
rect 2797 3484 2803 3536
rect 2733 3444 2739 3456
rect 2829 3424 2835 3556
rect 2893 3484 2899 3516
rect 2957 3484 2963 3676
rect 2973 3604 2979 3656
rect 2845 3477 2860 3483
rect 2845 3384 2851 3477
rect 2877 3464 2883 3476
rect 2941 3463 2947 3476
rect 2941 3457 2963 3463
rect 2957 3424 2963 3457
rect 2916 3417 2931 3423
rect 2861 3377 2899 3383
rect 2669 3304 2675 3356
rect 2797 3343 2803 3376
rect 2781 3337 2803 3343
rect 2708 3317 2723 3323
rect 2717 3304 2723 3317
rect 2701 3264 2707 3296
rect 2541 3177 2627 3183
rect 2637 3177 2659 3183
rect 2669 3237 2723 3243
rect 2461 3137 2483 3143
rect 2477 3084 2483 3137
rect 2493 3123 2499 3177
rect 2637 3163 2643 3177
rect 2509 3157 2643 3163
rect 2509 3144 2515 3157
rect 2653 3144 2659 3156
rect 2541 3124 2547 3136
rect 2493 3117 2515 3123
rect 2461 3063 2467 3076
rect 2461 3057 2483 3063
rect 2301 2943 2307 2956
rect 2349 2944 2355 2996
rect 2301 2937 2323 2943
rect 2317 2924 2323 2937
rect 2365 2904 2371 2996
rect 2381 2904 2387 2916
rect 2333 2864 2339 2896
rect 2356 2877 2380 2883
rect 2269 2783 2275 2836
rect 2253 2777 2275 2783
rect 2253 2744 2259 2777
rect 2285 2724 2291 2816
rect 2317 2717 2332 2723
rect 2317 2684 2323 2717
rect 2221 2677 2243 2683
rect 2253 2677 2268 2683
rect 2148 2577 2163 2583
rect 2173 2564 2179 2576
rect 2157 2543 2163 2556
rect 2189 2543 2195 2556
rect 2157 2537 2195 2543
rect 2125 2524 2131 2536
rect 2029 2364 2035 2476
rect 2093 2444 2099 2496
rect 2077 2304 2083 2416
rect 2109 2404 2115 2516
rect 2125 2364 2131 2516
rect 2205 2324 2211 2636
rect 2221 2624 2227 2677
rect 2253 2663 2259 2677
rect 2237 2657 2259 2663
rect 2237 2644 2243 2657
rect 2301 2643 2307 2676
rect 2365 2663 2371 2716
rect 2285 2637 2307 2643
rect 2349 2657 2371 2663
rect 2285 2543 2291 2637
rect 2349 2623 2355 2657
rect 2413 2644 2419 3036
rect 2445 2863 2451 2916
rect 2461 2884 2467 2916
rect 2445 2857 2467 2863
rect 2429 2784 2435 2816
rect 2445 2724 2451 2776
rect 2308 2617 2355 2623
rect 2301 2597 2348 2603
rect 2301 2564 2307 2597
rect 2285 2537 2307 2543
rect 2285 2404 2291 2516
rect 2301 2504 2307 2537
rect 2333 2504 2339 2536
rect 2221 2324 2227 2336
rect 2157 2317 2172 2323
rect 2157 2304 2163 2317
rect 2173 2284 2179 2296
rect 2237 2284 2243 2316
rect 2269 2284 2275 2396
rect 2301 2324 2307 2496
rect 2381 2484 2387 2616
rect 2413 2544 2419 2576
rect 2429 2564 2435 2656
rect 2445 2564 2451 2696
rect 2461 2683 2467 2857
rect 2477 2784 2483 3057
rect 2509 2924 2515 3117
rect 2669 3123 2675 3237
rect 2701 3124 2707 3216
rect 2653 3117 2675 3123
rect 2525 3063 2531 3096
rect 2541 3084 2547 3116
rect 2525 3057 2563 3063
rect 2525 3004 2531 3036
rect 2541 2904 2547 3036
rect 2557 3004 2563 3057
rect 2573 3044 2579 3076
rect 2589 3024 2595 3116
rect 2612 3097 2643 3103
rect 2637 3044 2643 3097
rect 2605 3024 2611 3036
rect 2573 2944 2579 2976
rect 2621 2963 2627 3036
rect 2653 3024 2659 3117
rect 2685 3103 2691 3116
rect 2685 3097 2700 3103
rect 2669 3044 2675 3096
rect 2685 2984 2691 3076
rect 2717 3043 2723 3237
rect 2733 3184 2739 3236
rect 2749 3144 2755 3316
rect 2781 3303 2787 3337
rect 2765 3297 2787 3303
rect 2765 3203 2771 3297
rect 2829 3303 2835 3336
rect 2820 3297 2835 3303
rect 2861 3303 2867 3377
rect 2893 3363 2899 3377
rect 2893 3357 2915 3363
rect 2909 3324 2915 3357
rect 2925 3303 2931 3417
rect 2941 3344 2947 3416
rect 2957 3324 2963 3396
rect 2973 3384 2979 3436
rect 2989 3424 2995 3757
rect 3037 3704 3043 3896
rect 3149 3884 3155 4036
rect 3165 3884 3171 3916
rect 3181 3904 3187 4036
rect 3172 3877 3187 3883
rect 3053 3764 3059 3856
rect 3069 3824 3075 3836
rect 3112 3806 3113 3814
rect 3121 3806 3123 3814
rect 3131 3806 3133 3814
rect 3141 3806 3143 3814
rect 3151 3806 3160 3814
rect 3181 3804 3187 3877
rect 3085 3784 3091 3796
rect 3197 3783 3203 4096
rect 3245 4063 3251 4116
rect 3261 4084 3267 4116
rect 3245 4057 3267 4063
rect 3261 3923 3267 4057
rect 3277 4023 3283 4136
rect 3277 4017 3299 4023
rect 3293 3984 3299 4017
rect 3261 3917 3283 3923
rect 3277 3884 3283 3917
rect 3181 3777 3203 3783
rect 3085 3684 3091 3696
rect 3005 3584 3011 3656
rect 3069 3624 3075 3676
rect 3021 3484 3027 3556
rect 3037 3464 3043 3476
rect 2852 3297 2867 3303
rect 2893 3297 2931 3303
rect 2781 3224 2787 3236
rect 2765 3197 2787 3203
rect 2781 3104 2787 3197
rect 2733 3064 2739 3096
rect 2797 3084 2803 3236
rect 2717 3037 2739 3043
rect 2733 2964 2739 3037
rect 2749 2984 2755 2996
rect 2765 2964 2771 3076
rect 2813 3064 2819 3216
rect 2829 3124 2835 3256
rect 2605 2957 2627 2963
rect 2589 2923 2595 2956
rect 2573 2917 2595 2923
rect 2509 2864 2515 2896
rect 2493 2704 2499 2756
rect 2509 2724 2515 2836
rect 2541 2724 2547 2776
rect 2557 2744 2563 2876
rect 2573 2784 2579 2917
rect 2589 2744 2595 2816
rect 2573 2723 2579 2736
rect 2605 2724 2611 2957
rect 2781 2944 2787 2956
rect 2701 2937 2716 2943
rect 2621 2923 2627 2936
rect 2621 2917 2643 2923
rect 2557 2717 2579 2723
rect 2541 2704 2547 2716
rect 2557 2704 2563 2717
rect 2621 2703 2627 2896
rect 2637 2803 2643 2917
rect 2637 2797 2659 2803
rect 2653 2764 2659 2797
rect 2701 2764 2707 2937
rect 2813 2943 2819 2996
rect 2845 2984 2851 3256
rect 2861 3104 2867 3116
rect 2877 3084 2883 3236
rect 2893 3224 2899 3297
rect 2941 3224 2947 3316
rect 2861 3004 2867 3076
rect 2804 2937 2819 2943
rect 2717 2917 2748 2923
rect 2717 2784 2723 2917
rect 2765 2923 2771 2936
rect 2765 2917 2803 2923
rect 2797 2863 2803 2917
rect 2820 2917 2851 2923
rect 2845 2903 2851 2917
rect 2845 2897 2860 2903
rect 2877 2883 2883 3056
rect 2909 3024 2915 3216
rect 2957 3143 2963 3216
rect 2973 3164 2979 3216
rect 2957 3137 2979 3143
rect 2941 3102 2947 3136
rect 2973 3124 2979 3137
rect 2973 3044 2979 3116
rect 2989 3044 2995 3296
rect 3005 3244 3011 3296
rect 3037 3184 3043 3236
rect 3053 3223 3059 3436
rect 3069 3363 3075 3596
rect 3101 3504 3107 3556
rect 3101 3484 3107 3496
rect 3117 3464 3123 3616
rect 3133 3444 3139 3676
rect 3149 3464 3155 3656
rect 3165 3584 3171 3696
rect 3181 3604 3187 3777
rect 3213 3723 3219 3836
rect 3261 3784 3267 3836
rect 3309 3764 3315 4156
rect 3373 3943 3379 4076
rect 3389 4064 3395 4296
rect 3565 4284 3571 4296
rect 3581 4284 3587 4316
rect 3645 4304 3651 4316
rect 3421 4264 3427 4276
rect 3421 4164 3427 4216
rect 3437 4124 3443 4196
rect 3469 4124 3475 4216
rect 3556 4177 3571 4183
rect 3565 4164 3571 4177
rect 3469 4084 3475 4116
rect 3405 3957 3484 3963
rect 3373 3937 3395 3943
rect 3373 3904 3379 3916
rect 3325 3844 3331 3896
rect 3389 3884 3395 3937
rect 3405 3924 3411 3957
rect 3453 3937 3491 3943
rect 3453 3924 3459 3937
rect 3485 3923 3491 3937
rect 3508 3937 3523 3943
rect 3485 3917 3507 3923
rect 3405 3863 3411 3896
rect 3389 3857 3411 3863
rect 3293 3737 3308 3743
rect 3293 3724 3299 3737
rect 3204 3717 3228 3723
rect 3261 3684 3267 3716
rect 3309 3704 3315 3716
rect 3325 3664 3331 3776
rect 3341 3724 3347 3836
rect 3389 3784 3395 3857
rect 3325 3584 3331 3596
rect 3213 3523 3219 3536
rect 3213 3517 3235 3523
rect 3172 3477 3187 3483
rect 3181 3424 3187 3477
rect 3229 3464 3235 3517
rect 3245 3483 3251 3556
rect 3245 3477 3260 3483
rect 3085 3383 3091 3416
rect 3112 3406 3113 3414
rect 3121 3406 3123 3414
rect 3131 3406 3133 3414
rect 3141 3406 3143 3414
rect 3151 3406 3160 3414
rect 3085 3377 3132 3383
rect 3181 3383 3187 3396
rect 3229 3384 3235 3436
rect 3172 3377 3187 3383
rect 3069 3357 3091 3363
rect 3085 3324 3091 3357
rect 3101 3304 3107 3336
rect 3053 3217 3091 3223
rect 3085 3184 3091 3217
rect 3076 3137 3091 3143
rect 3053 3063 3059 3136
rect 3085 3104 3091 3137
rect 3101 3084 3107 3176
rect 3149 3144 3155 3376
rect 3245 3323 3251 3477
rect 3261 3344 3267 3376
rect 3245 3317 3267 3323
rect 3117 3063 3123 3096
rect 3133 3084 3139 3116
rect 3053 3057 3123 3063
rect 3133 3057 3148 3063
rect 3133 3043 3139 3057
rect 3165 3044 3171 3316
rect 3236 3297 3244 3303
rect 3085 3037 3139 3043
rect 2941 2964 2947 3016
rect 3005 2984 3011 2996
rect 3069 2964 3075 3036
rect 2893 2957 2908 2963
rect 2893 2944 2899 2957
rect 2861 2877 2883 2883
rect 2797 2857 2851 2863
rect 2685 2723 2691 2756
rect 2669 2717 2691 2723
rect 2653 2704 2659 2716
rect 2621 2697 2643 2703
rect 2461 2677 2483 2683
rect 2461 2544 2467 2656
rect 2477 2603 2483 2677
rect 2500 2677 2508 2683
rect 2525 2683 2531 2696
rect 2525 2677 2540 2683
rect 2589 2677 2620 2683
rect 2557 2664 2563 2676
rect 2477 2597 2499 2603
rect 2493 2544 2499 2597
rect 2397 2524 2403 2536
rect 2397 2484 2403 2496
rect 2413 2484 2419 2536
rect 2365 2364 2371 2436
rect 2157 2224 2163 2276
rect 2333 2264 2339 2316
rect 2173 2243 2179 2256
rect 2269 2243 2275 2256
rect 2173 2237 2275 2243
rect 2189 2217 2227 2223
rect 2189 2204 2195 2217
rect 2221 2203 2227 2217
rect 2221 2197 2268 2203
rect 2013 2123 2019 2136
rect 2045 2124 2051 2176
rect 2013 2117 2028 2123
rect 2004 2097 2012 2103
rect 1997 1944 2003 2076
rect 1988 1917 2003 1923
rect 1789 1757 1827 1763
rect 1773 1737 1795 1743
rect 1741 1504 1747 1656
rect 1757 1584 1763 1596
rect 1677 1444 1683 1476
rect 1741 1464 1747 1476
rect 1613 1384 1619 1396
rect 1725 1384 1731 1456
rect 1741 1424 1747 1456
rect 1613 1304 1619 1336
rect 1661 1324 1667 1356
rect 1576 1206 1577 1214
rect 1585 1206 1587 1214
rect 1595 1206 1597 1214
rect 1605 1206 1607 1214
rect 1615 1206 1624 1214
rect 1549 1124 1555 1196
rect 1645 1124 1651 1256
rect 1725 1184 1731 1296
rect 1700 1157 1715 1163
rect 1709 1144 1715 1157
rect 1485 1023 1491 1096
rect 1549 1084 1555 1116
rect 1741 1104 1747 1396
rect 1757 1324 1763 1536
rect 1773 1484 1779 1516
rect 1789 1344 1795 1737
rect 1805 1704 1811 1716
rect 1821 1684 1827 1757
rect 1885 1743 1891 1856
rect 1901 1843 1907 1856
rect 1949 1844 1955 1896
rect 1997 1863 2003 1917
rect 2013 1883 2019 1936
rect 2061 1904 2067 2196
rect 2093 1903 2099 2156
rect 2109 2104 2115 2196
rect 2205 2157 2236 2163
rect 2157 2143 2163 2156
rect 2157 2137 2179 2143
rect 2141 1984 2147 2136
rect 2157 2104 2163 2137
rect 2173 2104 2179 2137
rect 2189 1984 2195 2136
rect 2205 2104 2211 2157
rect 2221 2004 2227 2136
rect 2253 2117 2268 2123
rect 2237 2104 2243 2116
rect 2253 2063 2259 2117
rect 2333 2123 2339 2156
rect 2365 2143 2371 2336
rect 2397 2184 2403 2376
rect 2413 2304 2419 2356
rect 2429 2344 2435 2496
rect 2413 2184 2419 2196
rect 2356 2137 2371 2143
rect 2333 2117 2355 2123
rect 2253 2057 2275 2063
rect 2269 2023 2275 2057
rect 2269 2017 2307 2023
rect 2301 1984 2307 2017
rect 2317 1983 2323 2116
rect 2333 2024 2339 2096
rect 2349 2024 2355 2117
rect 2365 2044 2371 2116
rect 2317 1977 2339 1983
rect 2077 1897 2099 1903
rect 2013 1877 2028 1883
rect 1997 1857 2035 1863
rect 1901 1837 1923 1843
rect 1869 1737 1891 1743
rect 1853 1643 1859 1736
rect 1869 1663 1875 1737
rect 1892 1717 1900 1723
rect 1917 1704 1923 1837
rect 1981 1784 1987 1836
rect 1997 1763 2003 1836
rect 2013 1784 2019 1816
rect 2029 1804 2035 1857
rect 2045 1844 2051 1896
rect 2077 1863 2083 1897
rect 2077 1857 2099 1863
rect 2045 1764 2051 1796
rect 2077 1784 2083 1836
rect 1997 1757 2028 1763
rect 1933 1704 1939 1756
rect 1965 1717 1980 1723
rect 1869 1657 1884 1663
rect 1853 1637 1891 1643
rect 1805 1623 1811 1636
rect 1805 1617 1827 1623
rect 1805 1504 1811 1536
rect 1821 1524 1827 1617
rect 1837 1617 1875 1623
rect 1837 1504 1843 1617
rect 1869 1583 1875 1617
rect 1885 1603 1891 1637
rect 1933 1604 1939 1656
rect 1885 1597 1923 1603
rect 1869 1577 1891 1583
rect 1885 1563 1891 1577
rect 1885 1557 1907 1563
rect 1901 1464 1907 1557
rect 1917 1464 1923 1597
rect 1949 1483 1955 1716
rect 1965 1684 1971 1717
rect 1965 1524 1971 1656
rect 1981 1584 1987 1696
rect 1997 1584 2003 1716
rect 1949 1477 1971 1483
rect 1805 1364 1811 1416
rect 1869 1364 1875 1456
rect 1949 1444 1955 1456
rect 1757 1124 1763 1236
rect 1789 1163 1795 1316
rect 1805 1184 1811 1356
rect 1885 1343 1891 1396
rect 1965 1384 1971 1477
rect 1981 1363 1987 1536
rect 2013 1524 2019 1696
rect 2029 1584 2035 1736
rect 2045 1604 2051 1716
rect 1997 1483 2003 1496
rect 1997 1477 2019 1483
rect 1949 1357 1987 1363
rect 1876 1337 1891 1343
rect 1789 1157 1811 1163
rect 1517 1024 1523 1076
rect 1469 1017 1491 1023
rect 1325 957 1363 963
rect 1325 803 1331 957
rect 1389 904 1395 996
rect 1469 964 1475 1017
rect 1453 944 1459 956
rect 1533 944 1539 1076
rect 1565 1024 1571 1056
rect 1597 964 1603 1016
rect 1613 924 1619 1076
rect 1645 984 1651 1076
rect 1677 1044 1683 1096
rect 1709 1084 1715 1096
rect 1789 1064 1795 1096
rect 1805 1084 1811 1157
rect 1821 1064 1827 1316
rect 1837 1184 1843 1276
rect 1853 1103 1859 1256
rect 1869 1184 1875 1196
rect 1885 1124 1891 1316
rect 1949 1284 1955 1357
rect 2013 1324 2019 1477
rect 2029 1423 2035 1476
rect 2045 1464 2051 1496
rect 2061 1484 2067 1776
rect 2093 1704 2099 1857
rect 2125 1744 2131 1956
rect 2173 1943 2179 1976
rect 2221 1943 2227 1956
rect 2173 1937 2227 1943
rect 2141 1904 2147 1916
rect 2157 1904 2163 1936
rect 2237 1924 2243 1936
rect 2180 1917 2211 1923
rect 2205 1903 2211 1917
rect 2253 1904 2259 1956
rect 2333 1944 2339 1977
rect 2205 1897 2236 1903
rect 2205 1883 2211 1897
rect 2317 1884 2323 1936
rect 2349 1924 2355 1976
rect 2381 1943 2387 2016
rect 2397 1984 2403 2016
rect 2429 1963 2435 2316
rect 2445 2264 2451 2436
rect 2477 2384 2483 2536
rect 2509 2523 2515 2636
rect 2493 2517 2515 2523
rect 2461 2204 2467 2336
rect 2493 2324 2499 2517
rect 2525 2384 2531 2636
rect 2589 2564 2595 2677
rect 2637 2664 2643 2697
rect 2605 2544 2611 2656
rect 2653 2624 2659 2676
rect 2621 2584 2627 2596
rect 2493 2184 2499 2276
rect 2445 1984 2451 2176
rect 2509 2163 2515 2376
rect 2557 2344 2563 2536
rect 2573 2324 2579 2536
rect 2637 2524 2643 2616
rect 2669 2563 2675 2717
rect 2749 2704 2755 2816
rect 2797 2744 2803 2836
rect 2765 2704 2771 2716
rect 2685 2584 2691 2656
rect 2749 2644 2755 2676
rect 2701 2604 2707 2636
rect 2669 2557 2691 2563
rect 2621 2384 2627 2496
rect 2525 2264 2531 2316
rect 2589 2304 2595 2336
rect 2605 2304 2611 2376
rect 2653 2364 2659 2536
rect 2669 2323 2675 2376
rect 2685 2344 2691 2557
rect 2701 2544 2707 2596
rect 2717 2544 2723 2556
rect 2765 2524 2771 2536
rect 2669 2317 2691 2323
rect 2573 2277 2588 2283
rect 2541 2263 2547 2276
rect 2573 2263 2579 2277
rect 2685 2264 2691 2317
rect 2541 2257 2579 2263
rect 2509 2157 2572 2163
rect 2621 2157 2652 2163
rect 2461 2124 2467 2156
rect 2493 2144 2499 2156
rect 2605 2144 2611 2156
rect 2541 2024 2547 2096
rect 2420 1957 2435 1963
rect 2365 1937 2387 1943
rect 2164 1877 2211 1883
rect 2269 1863 2275 1876
rect 2269 1857 2284 1863
rect 2292 1857 2307 1863
rect 2093 1604 2099 1676
rect 2093 1463 2099 1576
rect 2109 1524 2115 1656
rect 2125 1484 2131 1696
rect 2141 1544 2147 1816
rect 2157 1804 2163 1856
rect 2157 1704 2163 1756
rect 2173 1683 2179 1816
rect 2189 1784 2195 1816
rect 2157 1677 2179 1683
rect 2189 1757 2204 1763
rect 2157 1584 2163 1677
rect 2141 1484 2147 1516
rect 2125 1464 2131 1476
rect 2157 1464 2163 1496
rect 2093 1457 2115 1463
rect 2109 1423 2115 1457
rect 2029 1417 2051 1423
rect 2029 1364 2035 1396
rect 2029 1264 2035 1336
rect 1901 1104 1907 1236
rect 1917 1104 1923 1256
rect 2013 1123 2019 1236
rect 2045 1184 2051 1417
rect 2061 1417 2099 1423
rect 2109 1417 2131 1423
rect 2061 1284 2067 1417
rect 2093 1404 2099 1417
rect 2109 1344 2115 1356
rect 2125 1323 2131 1417
rect 2141 1364 2147 1456
rect 2173 1404 2179 1576
rect 2189 1504 2195 1757
rect 2253 1763 2259 1856
rect 2301 1823 2307 1857
rect 2333 1843 2339 1896
rect 2365 1884 2371 1937
rect 2381 1917 2451 1923
rect 2349 1863 2355 1876
rect 2349 1857 2364 1863
rect 2381 1844 2387 1917
rect 2445 1903 2451 1917
rect 2445 1897 2460 1903
rect 2333 1837 2355 1843
rect 2301 1817 2316 1823
rect 2349 1764 2355 1837
rect 2365 1764 2371 1796
rect 2397 1784 2403 1896
rect 2477 1884 2483 1976
rect 2253 1757 2275 1763
rect 2205 1664 2211 1736
rect 2237 1703 2243 1716
rect 2228 1697 2243 1703
rect 2221 1604 2227 1656
rect 2253 1623 2259 1736
rect 2237 1617 2259 1623
rect 2237 1584 2243 1617
rect 2269 1584 2275 1757
rect 2285 1757 2332 1763
rect 2285 1724 2291 1757
rect 2301 1683 2307 1736
rect 2317 1704 2323 1716
rect 2301 1677 2339 1683
rect 2285 1543 2291 1636
rect 2276 1537 2291 1543
rect 2301 1524 2307 1596
rect 2333 1524 2339 1677
rect 2349 1604 2355 1756
rect 2365 1723 2371 1756
rect 2381 1744 2387 1776
rect 2413 1744 2419 1836
rect 2429 1744 2435 1876
rect 2461 1863 2467 1876
rect 2461 1857 2476 1863
rect 2493 1803 2499 2016
rect 2573 1984 2579 2096
rect 2541 1944 2547 1976
rect 2589 1964 2595 2096
rect 2509 1823 2515 1876
rect 2541 1844 2547 1916
rect 2605 1864 2611 2036
rect 2621 2024 2627 2157
rect 2637 2044 2643 2136
rect 2685 2124 2691 2176
rect 2701 2144 2707 2516
rect 2717 2404 2723 2476
rect 2733 2384 2739 2516
rect 2781 2484 2787 2536
rect 2797 2524 2803 2576
rect 2797 2423 2803 2516
rect 2813 2444 2819 2756
rect 2845 2724 2851 2857
rect 2845 2564 2851 2656
rect 2861 2544 2867 2877
rect 2893 2864 2899 2896
rect 2877 2784 2883 2836
rect 2877 2584 2883 2616
rect 2893 2544 2899 2716
rect 2909 2704 2915 2916
rect 2925 2764 2931 2956
rect 2941 2924 2947 2956
rect 2941 2764 2947 2836
rect 2957 2784 2963 2916
rect 2973 2724 2979 2936
rect 2989 2924 2995 2956
rect 3005 2937 3020 2943
rect 3005 2903 3011 2937
rect 3044 2937 3075 2943
rect 2989 2897 3011 2903
rect 2989 2864 2995 2897
rect 3021 2864 3027 2916
rect 3053 2904 3059 2916
rect 3069 2884 3075 2937
rect 2989 2844 2995 2856
rect 2941 2563 2947 2716
rect 2989 2703 2995 2836
rect 3037 2824 3043 2876
rect 3085 2863 3091 3037
rect 3112 3006 3113 3014
rect 3121 3006 3123 3014
rect 3131 3006 3133 3014
rect 3141 3006 3143 3014
rect 3151 3006 3160 3014
rect 3181 2964 3187 3076
rect 3197 2964 3203 3136
rect 3213 3044 3219 3256
rect 3229 3243 3235 3256
rect 3229 3237 3244 3243
rect 3261 3184 3267 3317
rect 3277 3304 3283 3316
rect 3293 3183 3299 3376
rect 3309 3323 3315 3556
rect 3341 3504 3347 3656
rect 3357 3564 3363 3716
rect 3389 3624 3395 3716
rect 3405 3703 3411 3736
rect 3405 3697 3427 3703
rect 3421 3683 3427 3697
rect 3421 3677 3443 3683
rect 3373 3464 3379 3616
rect 3357 3324 3363 3436
rect 3373 3364 3379 3436
rect 3405 3363 3411 3656
rect 3421 3484 3427 3616
rect 3437 3504 3443 3677
rect 3453 3624 3459 3896
rect 3469 3884 3475 3916
rect 3485 3684 3491 3896
rect 3501 3663 3507 3917
rect 3517 3744 3523 3937
rect 3533 3924 3539 3936
rect 3549 3904 3555 3996
rect 3565 3944 3571 4076
rect 3581 3944 3587 4256
rect 3629 4184 3635 4196
rect 3645 4184 3651 4236
rect 3661 4143 3667 4476
rect 3677 4344 3683 4476
rect 3949 4464 3955 4536
rect 4141 4524 4147 4536
rect 4205 4504 4211 4516
rect 4141 4484 4147 4496
rect 3693 4284 3699 4356
rect 3741 4204 3747 4236
rect 3757 4184 3763 4316
rect 3885 4304 3891 4316
rect 3901 4284 3907 4456
rect 4077 4324 4083 4436
rect 3773 4184 3779 4196
rect 3789 4184 3795 4216
rect 3965 4184 3971 4316
rect 3997 4284 4003 4316
rect 4061 4302 4067 4303
rect 3684 4157 3724 4163
rect 3661 4137 3683 4143
rect 3613 4124 3619 4136
rect 3597 4064 3603 4116
rect 3613 4004 3619 4096
rect 3597 3984 3603 3996
rect 3645 3984 3651 3996
rect 3661 3923 3667 4116
rect 3677 4083 3683 4137
rect 3693 4104 3699 4136
rect 3709 4104 3715 4116
rect 3821 4104 3827 4136
rect 3837 4104 3843 4116
rect 3917 4104 3923 4116
rect 3933 4104 3939 4136
rect 3981 4123 3987 4236
rect 3997 4184 4003 4236
rect 4061 4184 4067 4294
rect 4084 4277 4092 4283
rect 4013 4157 4051 4163
rect 4013 4143 4019 4157
rect 4045 4144 4051 4157
rect 3972 4117 3987 4123
rect 3997 4137 4019 4143
rect 3677 4077 3699 4083
rect 3693 3984 3699 4077
rect 3709 3944 3715 4036
rect 3757 3924 3763 4096
rect 3796 4077 3843 4083
rect 3837 4064 3843 4077
rect 3805 4037 3884 4043
rect 3805 3943 3811 4037
rect 3901 3984 3907 3996
rect 3949 3944 3955 4096
rect 3997 4083 4003 4137
rect 4029 4124 4035 4136
rect 4077 4124 4083 4216
rect 4125 4164 4131 4256
rect 4157 4124 4163 4276
rect 4189 4264 4195 4336
rect 4205 4304 4211 4316
rect 4221 4264 4227 4436
rect 4253 4284 4259 4516
rect 4333 4384 4339 4516
rect 4349 4464 4355 4536
rect 4541 4504 4547 4516
rect 4413 4403 4419 4436
rect 4397 4397 4419 4403
rect 4397 4304 4403 4397
rect 4429 4384 4435 4496
rect 4509 4424 4515 4476
rect 4573 4464 4579 4536
rect 4941 4524 4947 4536
rect 4733 4484 4739 4516
rect 4781 4484 4787 4496
rect 4861 4464 4867 4476
rect 4509 4324 4515 4416
rect 4509 4304 4515 4316
rect 4301 4284 4307 4296
rect 3988 4077 4003 4083
rect 4013 3964 4019 4116
rect 3796 3937 3811 3943
rect 3988 3937 4003 3943
rect 3661 3917 3699 3923
rect 3693 3904 3699 3917
rect 3757 3904 3763 3916
rect 3636 3897 3651 3903
rect 3485 3657 3507 3663
rect 3485 3584 3491 3657
rect 3533 3564 3539 3776
rect 3469 3504 3475 3556
rect 3389 3357 3411 3363
rect 3389 3324 3395 3357
rect 3421 3344 3427 3396
rect 3309 3317 3331 3323
rect 3277 3177 3299 3183
rect 3277 3123 3283 3177
rect 3261 3117 3283 3123
rect 3069 2857 3091 2863
rect 3012 2757 3027 2763
rect 3021 2724 3027 2757
rect 3037 2724 3043 2816
rect 3053 2744 3059 2856
rect 3069 2784 3075 2857
rect 3101 2823 3107 2916
rect 3117 2864 3123 2956
rect 3229 2944 3235 3016
rect 3261 3004 3267 3117
rect 3325 3104 3331 3317
rect 3341 3184 3347 3316
rect 3357 3283 3363 3296
rect 3357 3277 3379 3283
rect 3341 3063 3347 3136
rect 3316 3057 3347 3063
rect 3357 3043 3363 3236
rect 3373 3223 3379 3277
rect 3389 3244 3395 3296
rect 3373 3217 3395 3223
rect 3389 3184 3395 3217
rect 3389 3064 3395 3156
rect 3309 3037 3363 3043
rect 3309 2983 3315 3037
rect 3268 2977 3315 2983
rect 3309 2944 3315 2956
rect 3165 2903 3171 2916
rect 3165 2897 3203 2903
rect 3197 2884 3203 2897
rect 3181 2863 3187 2876
rect 3229 2863 3235 2916
rect 3181 2857 3235 2863
rect 3085 2817 3107 2823
rect 3085 2723 3091 2817
rect 3101 2724 3107 2776
rect 3069 2717 3091 2723
rect 2973 2697 2995 2703
rect 2957 2604 2963 2696
rect 2925 2557 2947 2563
rect 2925 2544 2931 2557
rect 2973 2543 2979 2697
rect 3069 2684 3075 2717
rect 3117 2704 3123 2836
rect 3133 2684 3139 2856
rect 3165 2784 3171 2816
rect 3149 2704 3155 2716
rect 3181 2684 3187 2796
rect 2989 2624 2995 2676
rect 3005 2603 3011 2676
rect 3101 2644 3107 2676
rect 3117 2644 3123 2676
rect 3149 2643 3155 2676
rect 3197 2643 3203 2736
rect 3149 2637 3203 2643
rect 3037 2604 3043 2636
rect 2989 2597 3011 2603
rect 2989 2544 2995 2597
rect 3053 2564 3059 2616
rect 3069 2564 3075 2596
rect 3012 2557 3027 2563
rect 2964 2537 2979 2543
rect 2829 2524 2835 2536
rect 2845 2504 2851 2536
rect 2861 2484 2867 2536
rect 2941 2524 2947 2536
rect 2916 2517 2931 2523
rect 2836 2457 2867 2463
rect 2829 2423 2835 2436
rect 2797 2417 2835 2423
rect 2829 2363 2835 2376
rect 2861 2363 2867 2457
rect 2877 2444 2883 2516
rect 2925 2503 2931 2517
rect 2925 2497 2947 2503
rect 2829 2357 2867 2363
rect 2717 2184 2723 2276
rect 2733 2224 2739 2276
rect 2749 2184 2755 2256
rect 2765 2204 2771 2316
rect 2797 2284 2803 2356
rect 2877 2284 2883 2296
rect 2893 2284 2899 2496
rect 2909 2284 2915 2476
rect 2765 2164 2771 2176
rect 2797 2164 2803 2216
rect 2813 2144 2819 2156
rect 2653 2104 2659 2116
rect 2733 2104 2739 2136
rect 2653 2024 2659 2096
rect 2717 2024 2723 2096
rect 2621 1984 2627 1996
rect 2717 1963 2723 1996
rect 2749 1964 2755 2136
rect 2781 2003 2787 2076
rect 2797 2024 2803 2096
rect 2813 2064 2819 2116
rect 2781 1997 2803 2003
rect 2717 1957 2739 1963
rect 2557 1823 2563 1836
rect 2509 1817 2563 1823
rect 2573 1804 2579 1836
rect 2468 1797 2499 1803
rect 2589 1764 2595 1796
rect 2365 1717 2387 1723
rect 2189 1404 2195 1476
rect 2237 1463 2243 1516
rect 2365 1504 2371 1596
rect 2381 1584 2387 1717
rect 2420 1697 2435 1703
rect 2429 1684 2435 1697
rect 2397 1563 2403 1656
rect 2381 1557 2403 1563
rect 2381 1504 2387 1557
rect 2397 1504 2403 1516
rect 2413 1504 2419 1656
rect 2445 1524 2451 1676
rect 2461 1504 2467 1736
rect 2477 1564 2483 1716
rect 2509 1544 2515 1736
rect 2509 1504 2515 1516
rect 2253 1484 2259 1496
rect 2285 1464 2291 1476
rect 2228 1457 2243 1463
rect 2301 1384 2307 1496
rect 2317 1364 2323 1476
rect 2333 1424 2339 1496
rect 2413 1477 2428 1483
rect 2109 1317 2131 1323
rect 1997 1117 2019 1123
rect 1853 1097 1875 1103
rect 1853 1064 1859 1076
rect 1725 1057 1740 1063
rect 1709 1024 1715 1056
rect 1677 964 1683 1016
rect 1725 964 1731 1057
rect 1629 924 1635 956
rect 1533 903 1539 916
rect 1524 897 1539 903
rect 1485 883 1491 896
rect 1485 877 1500 883
rect 1341 864 1347 876
rect 1325 797 1347 803
rect 1341 744 1347 797
rect 1277 684 1283 736
rect 1373 704 1379 816
rect 1389 784 1395 796
rect 1437 764 1443 836
rect 1469 804 1475 836
rect 1517 784 1523 876
rect 1533 764 1539 897
rect 1549 824 1555 876
rect 1576 806 1577 814
rect 1585 806 1587 814
rect 1595 806 1597 814
rect 1605 806 1607 814
rect 1615 806 1624 814
rect 1645 764 1651 956
rect 1741 944 1747 1036
rect 1773 1004 1779 1056
rect 1805 1043 1811 1056
rect 1805 1037 1836 1043
rect 1757 924 1763 996
rect 1773 944 1779 956
rect 1469 757 1507 763
rect 989 677 1011 683
rect 925 564 931 636
rect 989 624 995 677
rect 1124 677 1132 683
rect 1037 624 1043 676
rect 957 564 963 616
rect 1053 584 1059 676
rect 925 524 931 556
rect 941 504 947 516
rect 957 483 963 496
rect 916 477 963 483
rect 989 320 995 358
rect 1053 344 1059 436
rect 1085 424 1091 516
rect 1085 324 1091 376
rect 1101 324 1107 636
rect 1117 604 1123 676
rect 1133 584 1139 656
rect 1165 564 1171 656
rect 1245 643 1251 676
rect 1245 637 1260 643
rect 1277 603 1283 616
rect 1261 597 1283 603
rect 1389 603 1395 756
rect 1469 744 1475 757
rect 1501 743 1507 757
rect 1501 737 1539 743
rect 1533 703 1539 737
rect 1437 697 1475 703
rect 1533 697 1571 703
rect 1437 683 1443 697
rect 1469 684 1475 697
rect 1565 684 1571 697
rect 1428 677 1443 683
rect 1389 597 1411 603
rect 1261 584 1267 597
rect 1197 564 1203 576
rect 1325 544 1331 576
rect 1389 544 1395 576
rect 1405 544 1411 597
rect 1140 537 1148 543
rect 1149 504 1155 516
rect 1117 423 1123 496
rect 1165 463 1171 516
rect 1213 483 1219 536
rect 1373 524 1379 536
rect 1437 524 1443 576
rect 1453 524 1459 656
rect 1533 644 1539 676
rect 1485 544 1491 636
rect 1469 524 1475 536
rect 1501 524 1507 536
rect 1405 504 1411 516
rect 1453 504 1459 516
rect 1325 497 1340 503
rect 1277 483 1283 496
rect 1213 477 1283 483
rect 1165 457 1203 463
rect 1149 437 1187 443
rect 1149 423 1155 437
rect 1181 424 1187 437
rect 1117 417 1155 423
rect 1149 304 1155 376
rect 1165 284 1171 416
rect 1197 324 1203 457
rect 1277 423 1283 477
rect 1277 417 1299 423
rect 1229 384 1235 396
rect 1229 344 1235 376
rect 1181 283 1187 316
rect 1261 284 1267 336
rect 1181 277 1212 283
rect 861 144 867 156
rect 253 62 259 116
rect 573 64 579 136
rect 877 124 883 216
rect 973 184 979 216
rect 925 144 931 176
rect 989 164 995 256
rect 1053 124 1059 196
rect 1069 184 1075 276
rect 893 117 908 123
rect 637 44 643 100
rect 845 103 851 116
rect 893 103 899 117
rect 973 104 979 116
rect 1069 104 1075 136
rect 1117 124 1123 236
rect 1197 204 1203 236
rect 1293 204 1299 417
rect 1309 284 1315 316
rect 1325 284 1331 497
rect 1373 324 1379 436
rect 1405 404 1411 496
rect 1421 404 1427 436
rect 1389 317 1404 323
rect 1389 303 1395 317
rect 1357 297 1395 303
rect 1341 284 1347 296
rect 1357 263 1363 297
rect 1453 284 1459 336
rect 1485 303 1491 496
rect 1517 424 1523 536
rect 1533 524 1539 636
rect 1549 584 1555 676
rect 1581 524 1587 736
rect 1597 524 1603 756
rect 1661 684 1667 916
rect 1677 804 1683 836
rect 1693 744 1699 896
rect 1613 603 1619 676
rect 1661 644 1667 676
rect 1725 644 1731 716
rect 1741 664 1747 816
rect 1757 724 1763 896
rect 1757 644 1763 696
rect 1773 684 1779 936
rect 1789 923 1795 1036
rect 1789 917 1811 923
rect 1805 723 1811 917
rect 1821 904 1827 1016
rect 1837 944 1843 956
rect 1796 717 1811 723
rect 1821 723 1827 836
rect 1853 724 1859 1036
rect 1869 1003 1875 1097
rect 1885 1043 1891 1096
rect 1885 1037 1907 1043
rect 1901 1024 1907 1037
rect 1869 997 1907 1003
rect 1901 984 1907 997
rect 1949 964 1955 1096
rect 1965 1064 1971 1096
rect 1981 1024 1987 1096
rect 1997 1084 2003 1117
rect 2061 1104 2067 1216
rect 2077 1184 2083 1316
rect 2013 1084 2019 1096
rect 1997 1024 2003 1076
rect 2077 1064 2083 1076
rect 1917 903 1923 956
rect 1997 924 2003 996
rect 1940 917 1971 923
rect 1901 897 1923 903
rect 1885 744 1891 896
rect 1821 717 1843 723
rect 1661 603 1667 616
rect 1613 597 1667 603
rect 1709 603 1715 636
rect 1709 597 1731 603
rect 1725 584 1731 597
rect 1581 444 1587 516
rect 1485 297 1500 303
rect 1517 284 1523 336
rect 1549 304 1555 436
rect 1576 406 1577 414
rect 1585 406 1587 414
rect 1595 406 1597 414
rect 1605 406 1607 414
rect 1615 406 1624 414
rect 1645 404 1651 536
rect 1661 523 1667 576
rect 1709 557 1747 563
rect 1684 537 1692 543
rect 1661 517 1699 523
rect 1613 357 1667 363
rect 1492 277 1500 283
rect 1533 283 1539 296
rect 1565 283 1571 296
rect 1533 277 1571 283
rect 1389 264 1395 276
rect 1341 257 1363 263
rect 1341 204 1347 257
rect 1437 244 1443 256
rect 1581 244 1587 356
rect 1597 244 1603 336
rect 1613 284 1619 357
rect 1661 324 1667 357
rect 1693 323 1699 517
rect 1709 504 1715 557
rect 1741 544 1747 557
rect 1725 524 1731 536
rect 1805 524 1811 676
rect 1821 623 1827 696
rect 1837 683 1843 717
rect 1869 683 1875 696
rect 1837 677 1875 683
rect 1821 617 1852 623
rect 1885 604 1891 636
rect 1901 583 1907 897
rect 1933 864 1939 896
rect 1949 864 1955 876
rect 1965 843 1971 917
rect 2013 883 2019 1056
rect 2061 1044 2067 1056
rect 1949 837 1971 843
rect 1997 877 2019 883
rect 1917 684 1923 796
rect 1933 744 1939 836
rect 1949 764 1955 837
rect 1997 744 2003 877
rect 2045 864 2051 976
rect 2061 964 2067 1016
rect 2077 1003 2083 1056
rect 2093 1024 2099 1316
rect 2109 1244 2115 1317
rect 2141 1144 2147 1356
rect 2237 1343 2243 1356
rect 2301 1344 2307 1356
rect 2237 1337 2300 1343
rect 2349 1343 2355 1416
rect 2333 1337 2355 1343
rect 2157 1324 2163 1336
rect 2157 1123 2163 1316
rect 2173 1304 2179 1316
rect 2173 1124 2179 1176
rect 2189 1143 2195 1316
rect 2221 1224 2227 1336
rect 2189 1137 2227 1143
rect 2141 1117 2163 1123
rect 2125 1104 2131 1116
rect 2141 1083 2147 1117
rect 2221 1123 2227 1137
rect 2221 1117 2243 1123
rect 2125 1077 2147 1083
rect 2077 997 2099 1003
rect 2093 943 2099 997
rect 2125 964 2131 1077
rect 2157 964 2163 1016
rect 2173 944 2179 1096
rect 2221 1084 2227 1096
rect 2189 1043 2195 1056
rect 2189 1037 2211 1043
rect 2068 937 2099 943
rect 2020 857 2028 863
rect 2029 704 2035 716
rect 1885 577 1907 583
rect 1869 544 1875 556
rect 1885 523 1891 577
rect 1901 524 1907 536
rect 1869 517 1891 523
rect 1853 504 1859 516
rect 1709 403 1715 436
rect 1741 404 1747 436
rect 1709 397 1731 403
rect 1725 324 1731 397
rect 1837 384 1843 496
rect 1796 337 1820 343
rect 1853 324 1859 436
rect 1869 404 1875 517
rect 1917 504 1923 676
rect 1933 624 1939 696
rect 2045 684 2051 816
rect 1949 524 1955 656
rect 1965 624 1971 636
rect 1981 604 1987 676
rect 2045 624 2051 636
rect 1965 544 1971 596
rect 2061 564 2067 736
rect 2093 723 2099 836
rect 2125 824 2131 856
rect 2141 824 2147 936
rect 2077 717 2099 723
rect 2077 704 2083 717
rect 2157 704 2163 716
rect 2173 704 2179 756
rect 2189 724 2195 1016
rect 2205 924 2211 1037
rect 2221 944 2227 1056
rect 2237 1023 2243 1117
rect 2253 1084 2259 1216
rect 2269 1084 2275 1236
rect 2301 1103 2307 1176
rect 2292 1097 2307 1103
rect 2317 1084 2323 1336
rect 2237 1017 2259 1023
rect 2253 1004 2259 1017
rect 2237 924 2243 996
rect 2269 964 2275 1056
rect 2333 1044 2339 1337
rect 2365 1244 2371 1396
rect 2397 1384 2403 1476
rect 2381 1324 2387 1356
rect 2397 1344 2403 1376
rect 2365 1163 2371 1216
rect 2381 1184 2387 1196
rect 2397 1163 2403 1316
rect 2413 1244 2419 1477
rect 2525 1483 2531 1756
rect 2509 1477 2531 1483
rect 2429 1424 2435 1456
rect 2445 1264 2451 1416
rect 2493 1344 2499 1456
rect 2509 1424 2515 1477
rect 2541 1443 2547 1756
rect 2605 1743 2611 1856
rect 2621 1763 2627 1916
rect 2637 1904 2643 1916
rect 2637 1884 2643 1896
rect 2653 1823 2659 1836
rect 2685 1823 2691 1916
rect 2701 1864 2707 1896
rect 2717 1884 2723 1936
rect 2733 1884 2739 1957
rect 2797 1924 2803 1997
rect 2813 1984 2819 2016
rect 2829 1963 2835 2256
rect 2845 2243 2851 2276
rect 2925 2264 2931 2376
rect 2941 2344 2947 2497
rect 2973 2444 2979 2537
rect 3021 2503 3027 2557
rect 3085 2523 3091 2616
rect 3112 2606 3113 2614
rect 3121 2606 3123 2614
rect 3131 2606 3133 2614
rect 3141 2606 3143 2614
rect 3151 2606 3160 2614
rect 3181 2564 3187 2616
rect 3197 2584 3203 2596
rect 3085 2517 3123 2523
rect 3005 2497 3027 2503
rect 2957 2324 2963 2416
rect 2989 2384 2995 2436
rect 3005 2304 3011 2497
rect 3069 2463 3075 2516
rect 3117 2503 3123 2517
rect 3117 2497 3139 2503
rect 3101 2464 3107 2496
rect 3133 2484 3139 2497
rect 3069 2457 3091 2463
rect 2893 2257 2908 2263
rect 2845 2237 2883 2243
rect 2877 2184 2883 2237
rect 2893 2184 2899 2257
rect 2941 2224 2947 2236
rect 2925 2163 2931 2216
rect 2973 2163 2979 2216
rect 2989 2163 2995 2296
rect 3005 2224 3011 2276
rect 3021 2264 3027 2416
rect 3037 2284 3043 2436
rect 3028 2237 3043 2243
rect 2925 2157 2963 2163
rect 2973 2157 2995 2163
rect 2845 1984 2851 2156
rect 2877 2144 2883 2156
rect 2925 2137 2940 2143
rect 2861 2084 2867 2116
rect 2861 1964 2867 2056
rect 2877 2024 2883 2056
rect 2893 2024 2899 2096
rect 2893 1964 2899 2016
rect 2829 1957 2851 1963
rect 2781 1864 2787 1896
rect 2813 1884 2819 1896
rect 2653 1817 2691 1823
rect 2621 1757 2636 1763
rect 2605 1737 2627 1743
rect 2621 1723 2627 1737
rect 2621 1717 2643 1723
rect 2605 1703 2611 1716
rect 2557 1697 2611 1703
rect 2557 1684 2563 1697
rect 2621 1684 2627 1696
rect 2589 1624 2595 1676
rect 2605 1663 2611 1676
rect 2605 1657 2627 1663
rect 2605 1624 2611 1636
rect 2589 1604 2595 1616
rect 2589 1544 2595 1556
rect 2525 1437 2547 1443
rect 2525 1363 2531 1437
rect 2509 1357 2531 1363
rect 2461 1283 2467 1296
rect 2461 1277 2483 1283
rect 2429 1204 2435 1236
rect 2365 1157 2403 1163
rect 2365 1084 2371 1116
rect 2381 1044 2387 1157
rect 2445 1124 2451 1236
rect 2477 1224 2483 1277
rect 2461 1123 2467 1136
rect 2461 1117 2483 1123
rect 2301 1037 2316 1043
rect 2205 764 2211 896
rect 2221 743 2227 916
rect 2237 764 2243 836
rect 2221 737 2243 743
rect 2205 723 2211 736
rect 2205 717 2227 723
rect 2189 703 2195 716
rect 2189 697 2204 703
rect 2093 684 2099 696
rect 2109 664 2115 676
rect 2109 644 2115 656
rect 2125 604 2131 696
rect 2221 684 2227 717
rect 2237 684 2243 737
rect 2253 703 2259 876
rect 2269 724 2275 916
rect 2285 824 2291 896
rect 2253 697 2268 703
rect 2285 703 2291 796
rect 2301 764 2307 1037
rect 2397 1024 2403 1116
rect 2413 1104 2419 1116
rect 2477 1104 2483 1117
rect 2404 997 2419 1003
rect 2333 944 2339 996
rect 2413 984 2419 997
rect 2429 964 2435 1056
rect 2461 1044 2467 1076
rect 2477 1064 2483 1096
rect 2493 1084 2499 1296
rect 2509 1284 2515 1357
rect 2557 1344 2563 1496
rect 2589 1464 2595 1496
rect 2589 1363 2595 1436
rect 2605 1424 2611 1516
rect 2621 1503 2627 1657
rect 2637 1544 2643 1717
rect 2717 1723 2723 1776
rect 2733 1743 2739 1816
rect 2733 1737 2755 1743
rect 2717 1717 2739 1723
rect 2669 1624 2675 1716
rect 2701 1664 2707 1716
rect 2733 1704 2739 1717
rect 2685 1603 2691 1616
rect 2669 1597 2691 1603
rect 2621 1497 2636 1503
rect 2589 1357 2611 1363
rect 2525 1304 2531 1336
rect 2557 1224 2563 1316
rect 2589 1304 2595 1336
rect 2605 1304 2611 1357
rect 2621 1324 2627 1497
rect 2653 1484 2659 1556
rect 2669 1504 2675 1597
rect 2701 1564 2707 1636
rect 2717 1624 2723 1696
rect 2749 1683 2755 1737
rect 2733 1677 2755 1683
rect 2733 1643 2739 1677
rect 2733 1637 2755 1643
rect 2692 1497 2707 1503
rect 2637 1443 2643 1476
rect 2637 1437 2659 1443
rect 2637 1364 2643 1376
rect 2653 1364 2659 1437
rect 2669 1424 2675 1436
rect 2701 1424 2707 1497
rect 2717 1383 2723 1476
rect 2669 1377 2723 1383
rect 2669 1344 2675 1377
rect 2653 1304 2659 1336
rect 2589 1284 2595 1296
rect 2685 1284 2691 1336
rect 2621 1263 2627 1276
rect 2621 1257 2643 1263
rect 2541 1123 2547 1216
rect 2589 1144 2595 1236
rect 2541 1117 2556 1123
rect 2509 1084 2515 1116
rect 2525 1104 2531 1116
rect 2605 1104 2611 1236
rect 2637 1163 2643 1257
rect 2653 1184 2659 1276
rect 2637 1157 2652 1163
rect 2541 1097 2556 1103
rect 2541 1064 2547 1097
rect 2621 1084 2627 1136
rect 2669 1123 2675 1236
rect 2701 1164 2707 1336
rect 2717 1324 2723 1336
rect 2733 1184 2739 1316
rect 2749 1124 2755 1637
rect 2765 1524 2771 1756
rect 2797 1704 2803 1776
rect 2813 1703 2819 1836
rect 2845 1784 2851 1957
rect 2925 1904 2931 2137
rect 2957 2143 2963 2157
rect 2957 2137 2979 2143
rect 2973 2124 2979 2137
rect 2989 2124 2995 2157
rect 2941 2084 2947 2116
rect 2957 2104 2963 2116
rect 3005 2104 3011 2136
rect 3037 2124 3043 2237
rect 3053 2184 3059 2356
rect 3085 2344 3091 2457
rect 3117 2324 3123 2476
rect 3181 2404 3187 2536
rect 3197 2524 3203 2576
rect 3213 2483 3219 2776
rect 3229 2743 3235 2836
rect 3245 2824 3251 2896
rect 3261 2844 3267 2936
rect 3277 2924 3283 2936
rect 3309 2803 3315 2936
rect 3341 2884 3347 3016
rect 3357 2964 3363 3016
rect 3405 2984 3411 3316
rect 3421 3264 3427 3316
rect 3437 3244 3443 3496
rect 3453 3484 3459 3496
rect 3533 3484 3539 3556
rect 3549 3484 3555 3876
rect 3581 3744 3587 3836
rect 3597 3723 3603 3836
rect 3613 3744 3619 3776
rect 3620 3737 3628 3743
rect 3645 3723 3651 3897
rect 3780 3897 3795 3903
rect 3725 3764 3731 3896
rect 3741 3783 3747 3896
rect 3773 3804 3779 3836
rect 3789 3784 3795 3897
rect 3741 3777 3763 3783
rect 3597 3717 3635 3723
rect 3613 3644 3619 3696
rect 3597 3484 3603 3636
rect 3629 3623 3635 3717
rect 3613 3617 3635 3623
rect 3645 3717 3660 3723
rect 3453 3364 3459 3456
rect 3469 3403 3475 3436
rect 3492 3417 3507 3423
rect 3469 3397 3491 3403
rect 3421 3164 3427 3236
rect 3453 3124 3459 3296
rect 3469 3264 3475 3376
rect 3485 3184 3491 3397
rect 3501 3383 3507 3417
rect 3517 3404 3523 3480
rect 3549 3464 3555 3476
rect 3613 3463 3619 3617
rect 3645 3543 3651 3717
rect 3629 3537 3651 3543
rect 3629 3484 3635 3537
rect 3661 3504 3667 3696
rect 3693 3524 3699 3536
rect 3709 3504 3715 3716
rect 3725 3683 3731 3736
rect 3741 3704 3747 3756
rect 3757 3683 3763 3777
rect 3725 3677 3763 3683
rect 3725 3524 3731 3556
rect 3613 3457 3635 3463
rect 3597 3384 3603 3416
rect 3501 3377 3555 3383
rect 3549 3364 3555 3377
rect 3533 3344 3539 3356
rect 3501 3184 3507 3316
rect 3421 2963 3427 3116
rect 3444 3077 3459 3083
rect 3405 2957 3427 2963
rect 3357 2944 3363 2956
rect 3405 2924 3411 2957
rect 3437 2944 3443 3056
rect 3453 3044 3459 3077
rect 3469 2984 3475 3036
rect 3453 2944 3459 2976
rect 3469 2904 3475 2956
rect 3412 2897 3459 2903
rect 3389 2857 3443 2863
rect 3293 2797 3315 2803
rect 3293 2784 3299 2797
rect 3229 2737 3251 2743
rect 3245 2683 3251 2737
rect 3277 2737 3292 2743
rect 3261 2704 3267 2736
rect 3277 2704 3283 2737
rect 3245 2677 3267 2683
rect 3236 2637 3251 2643
rect 3245 2564 3251 2637
rect 3261 2603 3267 2677
rect 3277 2644 3283 2676
rect 3293 2644 3299 2716
rect 3309 2664 3315 2776
rect 3325 2724 3331 2836
rect 3357 2764 3363 2836
rect 3373 2823 3379 2856
rect 3389 2844 3395 2857
rect 3373 2817 3395 2823
rect 3332 2697 3356 2703
rect 3373 2684 3379 2756
rect 3389 2684 3395 2817
rect 3405 2784 3411 2836
rect 3437 2744 3443 2857
rect 3453 2844 3459 2897
rect 3485 2763 3491 3116
rect 3533 3104 3539 3316
rect 3549 3204 3555 3316
rect 3533 3084 3539 3096
rect 3581 3084 3587 3356
rect 3597 3303 3603 3336
rect 3613 3324 3619 3356
rect 3629 3344 3635 3457
rect 3677 3423 3683 3456
rect 3668 3417 3683 3423
rect 3693 3404 3699 3496
rect 3725 3464 3731 3496
rect 3716 3437 3731 3443
rect 3725 3424 3731 3437
rect 3741 3424 3747 3536
rect 3757 3464 3763 3496
rect 3773 3444 3779 3756
rect 3789 3584 3795 3756
rect 3821 3744 3827 3916
rect 3917 3897 3932 3903
rect 3805 3704 3811 3736
rect 3821 3704 3827 3716
rect 3821 3503 3827 3696
rect 3837 3684 3843 3836
rect 3853 3784 3859 3836
rect 3885 3804 3891 3856
rect 3853 3703 3859 3756
rect 3917 3724 3923 3897
rect 3949 3864 3955 3916
rect 3997 3903 4003 3937
rect 4013 3924 4019 3936
rect 4045 3923 4051 3996
rect 4077 3984 4083 4076
rect 4093 3944 4099 4076
rect 4157 3944 4163 4096
rect 4173 4084 4179 4096
rect 4068 3937 4076 3943
rect 4029 3917 4051 3923
rect 4029 3903 4035 3917
rect 4084 3917 4115 3923
rect 4109 3903 4115 3917
rect 3997 3897 4035 3903
rect 4061 3897 4099 3903
rect 4109 3897 4124 3903
rect 3981 3863 3987 3896
rect 4061 3884 4067 3897
rect 4093 3884 4099 3897
rect 3981 3857 4012 3863
rect 3997 3823 4003 3836
rect 3981 3817 4003 3823
rect 3981 3804 3987 3817
rect 3997 3724 4003 3796
rect 4077 3724 4083 3876
rect 4157 3864 4163 3876
rect 4173 3804 4179 3896
rect 4189 3864 4195 4236
rect 4269 4203 4275 4276
rect 4253 4197 4275 4203
rect 4237 4083 4243 4116
rect 4253 4104 4259 4197
rect 4285 4103 4291 4216
rect 4381 4164 4387 4296
rect 4397 4204 4403 4296
rect 4461 4263 4467 4276
rect 4445 4257 4467 4263
rect 4413 4177 4428 4183
rect 4413 4164 4419 4177
rect 4445 4144 4451 4257
rect 4317 4104 4323 4136
rect 4525 4124 4531 4236
rect 4541 4144 4547 4456
rect 4664 4406 4665 4414
rect 4673 4406 4675 4414
rect 4683 4406 4685 4414
rect 4693 4406 4695 4414
rect 4703 4406 4712 4414
rect 4589 4124 4595 4276
rect 4605 4224 4611 4296
rect 4653 4284 4659 4316
rect 4701 4304 4707 4316
rect 4957 4304 4963 4536
rect 5021 4444 5027 4516
rect 5053 4444 5059 4456
rect 5053 4304 5059 4436
rect 5117 4423 5123 4496
rect 5245 4464 5251 4536
rect 5357 4524 5363 4556
rect 5101 4417 5123 4423
rect 5101 4324 5107 4417
rect 4621 4184 4627 4236
rect 4685 4164 4691 4276
rect 4749 4244 4755 4276
rect 4861 4264 4867 4296
rect 4909 4284 4915 4296
rect 4813 4177 4828 4183
rect 4813 4164 4819 4177
rect 4957 4164 4963 4296
rect 5053 4284 5059 4296
rect 4717 4124 4723 4136
rect 5053 4124 5059 4176
rect 5101 4143 5107 4316
rect 5149 4223 5155 4416
rect 5373 4384 5379 4536
rect 5549 4524 5555 4536
rect 5613 4524 5619 4556
rect 5741 4524 5747 4536
rect 5412 4517 5420 4523
rect 5588 4517 5603 4523
rect 5597 4504 5603 4517
rect 5613 4504 5619 4516
rect 5757 4504 5763 4516
rect 5789 4504 5795 4516
rect 5165 4284 5171 4316
rect 5229 4304 5235 4356
rect 5389 4324 5395 4496
rect 5453 4484 5459 4496
rect 5469 4364 5475 4436
rect 5392 4317 5395 4324
rect 5469 4323 5475 4356
rect 5485 4344 5491 4496
rect 5501 4464 5507 4496
rect 5581 4464 5587 4496
rect 5677 4484 5683 4496
rect 5453 4317 5475 4323
rect 5453 4304 5459 4317
rect 5485 4303 5491 4336
rect 5549 4323 5555 4456
rect 5629 4444 5635 4476
rect 5709 4364 5715 4496
rect 5757 4484 5763 4496
rect 5789 4384 5795 4456
rect 5629 4324 5635 4336
rect 5757 4324 5763 4356
rect 5533 4317 5555 4323
rect 5517 4304 5523 4316
rect 5469 4297 5491 4303
rect 5181 4284 5187 4296
rect 5357 4284 5363 4296
rect 5373 4284 5379 4296
rect 5469 4284 5475 4297
rect 5533 4284 5539 4317
rect 5581 4284 5587 4296
rect 5245 4243 5251 4276
rect 5245 4237 5267 4243
rect 5133 4217 5155 4223
rect 5117 4144 5123 4156
rect 5092 4137 5107 4143
rect 4285 4097 4307 4103
rect 4301 4084 4307 4097
rect 4237 4077 4259 4083
rect 4221 4023 4227 4076
rect 4205 4017 4227 4023
rect 4205 3944 4211 4017
rect 4221 4004 4227 4017
rect 4253 3904 4259 4077
rect 4285 4004 4291 4076
rect 4349 4004 4355 4076
rect 4285 3904 4291 3976
rect 4349 3924 4355 3976
rect 4349 3884 4355 3896
rect 4157 3783 4163 3796
rect 4157 3777 4172 3783
rect 3853 3697 3875 3703
rect 3837 3584 3843 3596
rect 3812 3497 3827 3503
rect 3853 3464 3859 3496
rect 3661 3344 3667 3356
rect 3629 3303 3635 3336
rect 3677 3323 3683 3396
rect 3821 3384 3827 3456
rect 3869 3383 3875 3697
rect 3917 3544 3923 3716
rect 3933 3624 3939 3716
rect 3901 3483 3907 3516
rect 3917 3504 3923 3516
rect 3901 3477 3939 3483
rect 3853 3377 3875 3383
rect 3805 3344 3811 3356
rect 3757 3337 3772 3343
rect 3661 3317 3683 3323
rect 3597 3297 3619 3303
rect 3629 3297 3651 3303
rect 3613 3124 3619 3297
rect 3645 3104 3651 3297
rect 3661 3164 3667 3317
rect 3757 3323 3763 3337
rect 3748 3317 3763 3323
rect 3693 3303 3699 3316
rect 3693 3297 3724 3303
rect 3773 3303 3779 3316
rect 3821 3304 3827 3356
rect 3853 3324 3859 3377
rect 3885 3324 3891 3436
rect 3933 3423 3939 3477
rect 3949 3444 3955 3716
rect 3981 3704 3987 3716
rect 4093 3704 4099 3756
rect 4157 3704 4163 3716
rect 4173 3704 4179 3736
rect 4061 3684 4067 3696
rect 4125 3684 4131 3696
rect 4020 3677 4044 3683
rect 4013 3617 4051 3623
rect 4013 3603 4019 3617
rect 3965 3597 4019 3603
rect 3965 3564 3971 3597
rect 4045 3603 4051 3617
rect 4045 3597 4060 3603
rect 3981 3544 3987 3556
rect 3972 3517 4012 3523
rect 4029 3503 4035 3596
rect 4061 3544 4067 3556
rect 4093 3524 4099 3556
rect 4141 3544 4147 3636
rect 4173 3524 4179 3696
rect 4189 3684 4195 3796
rect 4333 3777 4348 3783
rect 4205 3703 4211 3736
rect 4237 3724 4243 3736
rect 4205 3697 4227 3703
rect 4221 3603 4227 3697
rect 4253 3684 4259 3776
rect 4333 3764 4339 3777
rect 4509 3744 4515 3876
rect 4589 3824 4595 4116
rect 4701 4064 4707 4116
rect 4941 4104 4947 4116
rect 4664 4006 4665 4014
rect 4673 4006 4675 4014
rect 4683 4006 4685 4014
rect 4693 4006 4695 4014
rect 4703 4006 4712 4014
rect 4637 3984 4643 3996
rect 4957 3902 4963 4116
rect 5021 3944 5027 4096
rect 5085 3944 5091 4136
rect 5053 3924 5059 3936
rect 5133 3924 5139 4217
rect 5181 4124 5187 4176
rect 5245 4144 5251 4196
rect 5261 4144 5267 4237
rect 5277 4184 5283 4236
rect 5341 4224 5347 4276
rect 5357 4203 5363 4276
rect 5565 4263 5571 4276
rect 5597 4263 5603 4276
rect 5613 4264 5619 4296
rect 5661 4284 5667 4296
rect 5693 4264 5699 4316
rect 5789 4304 5795 4336
rect 5821 4324 5827 4356
rect 5837 4324 5843 4496
rect 5869 4384 5875 4536
rect 5917 4524 5923 4577
rect 5933 4544 5939 4556
rect 5997 4544 6003 4556
rect 5885 4424 5891 4496
rect 5869 4363 5875 4376
rect 5949 4364 5955 4536
rect 5981 4484 5987 4496
rect 5997 4404 6003 4536
rect 6013 4524 6019 4556
rect 6045 4424 6051 4496
rect 6061 4444 6067 4516
rect 6093 4483 6099 4536
rect 6173 4524 6179 4576
rect 6109 4504 6115 4516
rect 6093 4477 6115 4483
rect 6029 4384 6035 4396
rect 5853 4357 5875 4363
rect 5853 4344 5859 4357
rect 5837 4317 5840 4324
rect 5757 4284 5763 4296
rect 5741 4264 5747 4276
rect 5565 4257 5603 4263
rect 5341 4197 5363 4203
rect 5341 4144 5347 4197
rect 5389 4184 5395 4216
rect 5229 4104 5235 4136
rect 5389 4124 5395 4176
rect 5485 4163 5491 4236
rect 5501 4224 5507 4256
rect 5549 4184 5555 4236
rect 5725 4184 5731 4256
rect 5485 4157 5507 4163
rect 5437 4124 5443 4156
rect 5485 4124 5491 4136
rect 5501 4124 5507 4157
rect 5661 4144 5667 4176
rect 5789 4144 5795 4256
rect 5805 4224 5811 4276
rect 5853 4244 5859 4296
rect 5869 4284 5875 4336
rect 5885 4324 5891 4336
rect 5917 4323 5923 4336
rect 5917 4317 5955 4323
rect 5901 4284 5907 4316
rect 5949 4304 5955 4317
rect 5684 4137 5692 4143
rect 5213 4064 5219 4096
rect 5181 4024 5187 4036
rect 4701 3824 4707 3856
rect 4557 3744 4563 3756
rect 4285 3724 4291 3736
rect 4221 3597 4259 3603
rect 4253 3564 4259 3597
rect 3972 3497 4076 3503
rect 3965 3423 3971 3436
rect 3981 3424 3987 3436
rect 3933 3417 3971 3423
rect 4029 3383 4035 3456
rect 4125 3444 4131 3496
rect 4205 3484 4211 3536
rect 4237 3524 4243 3556
rect 4237 3504 4243 3516
rect 4301 3504 4307 3716
rect 4381 3564 4387 3616
rect 4141 3423 4147 3436
rect 4125 3417 4147 3423
rect 4029 3377 4044 3383
rect 3773 3297 3795 3303
rect 3677 3184 3683 3296
rect 3693 3164 3699 3276
rect 3725 3263 3731 3296
rect 3725 3257 3779 3263
rect 3773 3244 3779 3257
rect 3677 3143 3683 3156
rect 3668 3137 3683 3143
rect 3741 3084 3747 3196
rect 3652 3077 3667 3083
rect 3533 2944 3539 3076
rect 3581 2984 3587 3036
rect 3597 2924 3603 2956
rect 3613 2904 3619 2936
rect 3645 2904 3651 3056
rect 3661 3004 3667 3077
rect 3716 3077 3740 3083
rect 3693 3004 3699 3076
rect 3757 3004 3763 3236
rect 3789 3144 3795 3297
rect 3773 3103 3779 3136
rect 3805 3104 3811 3236
rect 3837 3217 3875 3223
rect 3821 3124 3827 3136
rect 3773 3097 3795 3103
rect 3789 3083 3795 3097
rect 3837 3103 3843 3217
rect 3869 3204 3875 3217
rect 3853 3144 3859 3196
rect 3821 3097 3843 3103
rect 3821 3083 3827 3097
rect 3853 3084 3859 3136
rect 3933 3104 3939 3276
rect 3965 3244 3971 3316
rect 4077 3303 4083 3336
rect 4068 3297 4083 3303
rect 3965 3157 4003 3163
rect 3965 3143 3971 3157
rect 3997 3144 4003 3157
rect 4029 3144 4035 3296
rect 4093 3283 4099 3336
rect 4109 3304 4115 3336
rect 4093 3277 4115 3283
rect 4093 3164 4099 3236
rect 4109 3163 4115 3277
rect 4125 3204 4131 3417
rect 4141 3344 4147 3396
rect 4205 3384 4211 3396
rect 4157 3304 4163 3336
rect 4164 3297 4179 3303
rect 4173 3203 4179 3297
rect 4189 3223 4195 3336
rect 4269 3324 4275 3416
rect 4301 3384 4307 3496
rect 4333 3464 4339 3536
rect 4461 3444 4467 3496
rect 4477 3484 4483 3736
rect 4557 3724 4563 3736
rect 4621 3603 4627 3816
rect 4941 3784 4947 3876
rect 4909 3724 4915 3756
rect 4941 3744 4947 3776
rect 4973 3744 4979 3816
rect 4989 3784 4995 3916
rect 5053 3904 5059 3916
rect 5085 3744 5091 3796
rect 5101 3744 5107 3876
rect 5133 3804 5139 3916
rect 5197 3904 5203 3916
rect 5229 3884 5235 4096
rect 5245 3884 5251 3916
rect 5325 3884 5331 3916
rect 5373 3884 5379 3996
rect 5485 3904 5491 4056
rect 5517 3903 5523 4136
rect 5677 4104 5683 4116
rect 5741 4104 5747 4136
rect 5741 3924 5747 3936
rect 5613 3917 5628 3923
rect 5501 3897 5523 3903
rect 5405 3884 5411 3896
rect 5181 3864 5187 3876
rect 5373 3864 5379 3876
rect 5453 3864 5459 3896
rect 5501 3884 5507 3897
rect 5597 3884 5603 3896
rect 5533 3864 5539 3876
rect 5613 3864 5619 3917
rect 5636 3917 5660 3923
rect 5661 3884 5667 3896
rect 5197 3784 5203 3796
rect 5261 3784 5267 3816
rect 4829 3704 4835 3716
rect 4637 3637 4668 3643
rect 4637 3624 4643 3637
rect 4708 3637 4739 3643
rect 4664 3606 4665 3614
rect 4673 3606 4675 3614
rect 4683 3606 4685 3614
rect 4693 3606 4695 3614
rect 4703 3606 4712 3614
rect 4621 3597 4643 3603
rect 4589 3564 4595 3596
rect 4589 3504 4595 3516
rect 4637 3504 4643 3597
rect 4733 3583 4739 3637
rect 4724 3577 4739 3583
rect 4893 3524 4899 3536
rect 4333 3344 4339 3376
rect 4349 3344 4355 3376
rect 4477 3364 4483 3476
rect 4733 3464 4739 3516
rect 4845 3504 4851 3516
rect 4781 3464 4787 3476
rect 4557 3383 4563 3456
rect 4548 3377 4563 3383
rect 4477 3344 4483 3356
rect 4605 3324 4611 3336
rect 4621 3324 4627 3436
rect 4765 3384 4771 3456
rect 4749 3364 4755 3376
rect 4781 3363 4787 3456
rect 4765 3357 4787 3363
rect 4413 3317 4428 3323
rect 4269 3304 4275 3316
rect 4413 3304 4419 3317
rect 4189 3217 4211 3223
rect 4157 3197 4179 3203
rect 4205 3203 4211 3217
rect 4205 3197 4227 3203
rect 4141 3163 4147 3196
rect 4109 3157 4147 3163
rect 3949 3137 3971 3143
rect 3949 3104 3955 3137
rect 4125 3124 4131 3136
rect 4157 3124 4163 3197
rect 4221 3163 4227 3197
rect 4237 3184 4243 3216
rect 4333 3197 4403 3203
rect 4333 3163 4339 3197
rect 4397 3184 4403 3197
rect 4221 3157 4339 3163
rect 4173 3124 4179 3136
rect 4429 3124 4435 3296
rect 4388 3117 4403 3123
rect 4084 3097 4099 3103
rect 3869 3084 3875 3096
rect 3933 3084 3939 3096
rect 3789 3077 3827 3083
rect 3892 3077 3907 3083
rect 3773 3064 3779 3076
rect 3837 3057 3875 3063
rect 3693 2977 3756 2983
rect 3677 2944 3683 2956
rect 3693 2944 3699 2977
rect 3661 2904 3667 2916
rect 3549 2864 3555 2896
rect 3517 2784 3523 2796
rect 3565 2764 3571 2796
rect 3581 2784 3587 2816
rect 3597 2764 3603 2896
rect 3469 2757 3491 2763
rect 3261 2597 3283 2603
rect 3261 2564 3267 2576
rect 3197 2477 3219 2483
rect 3197 2404 3203 2477
rect 3101 2244 3107 2296
rect 3117 2264 3123 2296
rect 3213 2244 3219 2456
rect 3229 2424 3235 2476
rect 3229 2264 3235 2376
rect 3021 2103 3027 2116
rect 3021 2097 3043 2103
rect 2989 2064 2995 2096
rect 2893 1803 2899 1876
rect 2973 1844 2979 2016
rect 3021 1984 3027 2076
rect 3037 2064 3043 2097
rect 3069 1984 3075 2156
rect 3085 2144 3091 2216
rect 3112 2206 3113 2214
rect 3121 2206 3123 2214
rect 3131 2206 3133 2214
rect 3141 2206 3143 2214
rect 3151 2206 3160 2214
rect 3101 1984 3107 2176
rect 3101 1924 3107 1956
rect 3117 1924 3123 2136
rect 3181 2124 3187 2196
rect 3213 2184 3219 2216
rect 3229 2163 3235 2256
rect 3213 2157 3235 2163
rect 3213 2123 3219 2157
rect 3213 2117 3235 2123
rect 3133 2023 3139 2096
rect 3149 2023 3155 2096
rect 3165 2084 3171 2116
rect 3133 2017 3155 2023
rect 3133 1983 3139 2017
rect 3149 1983 3155 2017
rect 3181 1984 3187 2016
rect 3133 1977 3155 1983
rect 2989 1823 2995 1896
rect 2884 1797 2899 1803
rect 2973 1817 2995 1823
rect 2973 1784 2979 1817
rect 3085 1784 3091 1896
rect 3149 1884 3155 1977
rect 3197 1904 3203 2016
rect 3213 1984 3219 2096
rect 3181 1883 3187 1896
rect 3181 1877 3203 1883
rect 3112 1806 3113 1814
rect 3121 1806 3123 1814
rect 3131 1806 3133 1814
rect 3141 1806 3143 1814
rect 3151 1806 3160 1814
rect 2989 1764 2995 1776
rect 2829 1724 2835 1736
rect 2877 1724 2883 1756
rect 2813 1697 2835 1703
rect 2781 1603 2787 1696
rect 2829 1624 2835 1697
rect 2845 1684 2851 1696
rect 2861 1624 2867 1696
rect 2893 1664 2899 1696
rect 2925 1643 2931 1736
rect 2973 1704 2979 1756
rect 2909 1637 2931 1643
rect 2781 1597 2803 1603
rect 2797 1583 2803 1597
rect 2861 1584 2867 1596
rect 2797 1577 2835 1583
rect 2781 1537 2819 1543
rect 2781 1504 2787 1537
rect 2797 1504 2803 1516
rect 2813 1504 2819 1537
rect 2829 1484 2835 1577
rect 2765 1384 2771 1416
rect 2781 1344 2787 1376
rect 2813 1344 2819 1476
rect 2829 1364 2835 1456
rect 2845 1344 2851 1516
rect 2861 1384 2867 1476
rect 2877 1424 2883 1496
rect 2893 1484 2899 1496
rect 2861 1344 2867 1376
rect 2772 1317 2780 1323
rect 2669 1117 2707 1123
rect 2564 1057 2627 1063
rect 2621 1044 2627 1057
rect 2644 1057 2691 1063
rect 2477 1023 2483 1036
rect 2461 1017 2483 1023
rect 2461 964 2467 1017
rect 2525 997 2595 1003
rect 2445 957 2460 963
rect 2356 917 2371 923
rect 2317 724 2323 876
rect 2340 817 2355 823
rect 2320 717 2323 724
rect 2285 697 2307 703
rect 2180 677 2211 683
rect 2173 644 2179 656
rect 2189 623 2195 636
rect 2141 617 2195 623
rect 2205 623 2211 677
rect 2253 677 2284 683
rect 2221 663 2227 676
rect 2253 663 2259 677
rect 2221 657 2259 663
rect 2205 617 2259 623
rect 1997 524 2003 556
rect 2036 517 2051 523
rect 1885 324 1891 396
rect 1693 317 1715 323
rect 1629 284 1635 316
rect 1677 303 1683 316
rect 1661 297 1683 303
rect 1661 263 1667 297
rect 1709 284 1715 317
rect 1869 304 1875 316
rect 1732 297 1756 303
rect 1773 297 1836 303
rect 1773 283 1779 297
rect 1901 284 1907 296
rect 1917 284 1923 496
rect 1981 464 1987 496
rect 2045 483 2051 517
rect 2045 477 2067 483
rect 2013 464 2019 476
rect 2061 464 2067 477
rect 1933 343 1939 456
rect 1933 337 1955 343
rect 1933 304 1939 316
rect 1949 304 1955 337
rect 1972 337 2003 343
rect 1997 304 2003 337
rect 2093 304 2099 556
rect 2109 544 2115 596
rect 2125 524 2131 576
rect 2141 504 2147 617
rect 2157 523 2163 556
rect 2189 524 2195 556
rect 2205 524 2211 536
rect 2157 517 2179 523
rect 2173 503 2179 517
rect 2221 504 2227 536
rect 2237 524 2243 596
rect 2253 563 2259 617
rect 2253 557 2268 563
rect 2301 524 2307 697
rect 2333 664 2339 716
rect 2349 544 2355 817
rect 2365 584 2371 917
rect 2381 864 2387 956
rect 2397 704 2403 836
rect 2413 703 2419 956
rect 2445 744 2451 957
rect 2468 937 2492 943
rect 2525 923 2531 997
rect 2589 983 2595 997
rect 2589 977 2611 983
rect 2605 964 2611 977
rect 2541 943 2547 956
rect 2589 944 2595 956
rect 2541 937 2579 943
rect 2525 917 2540 923
rect 2477 764 2483 836
rect 2493 764 2499 916
rect 2525 904 2531 917
rect 2573 923 2579 937
rect 2573 917 2595 923
rect 2589 904 2595 917
rect 2548 897 2563 903
rect 2557 883 2563 897
rect 2653 883 2659 956
rect 2557 877 2579 883
rect 2461 724 2467 736
rect 2413 697 2460 703
rect 2493 703 2499 756
rect 2525 704 2531 736
rect 2493 697 2508 703
rect 2381 564 2387 636
rect 2317 524 2323 536
rect 2285 504 2291 516
rect 2173 497 2211 503
rect 2205 483 2211 497
rect 2333 503 2339 536
rect 2365 524 2371 556
rect 2397 544 2403 676
rect 2445 584 2451 676
rect 2493 563 2499 676
rect 2541 663 2547 776
rect 2557 684 2563 856
rect 2573 744 2579 877
rect 2637 877 2659 883
rect 2589 704 2595 716
rect 2573 683 2579 696
rect 2573 677 2595 683
rect 2525 657 2547 663
rect 2525 644 2531 657
rect 2493 557 2515 563
rect 2445 543 2451 556
rect 2445 537 2467 543
rect 2429 503 2435 516
rect 2333 497 2435 503
rect 2205 477 2227 483
rect 2221 464 2227 477
rect 2205 443 2211 456
rect 2205 437 2275 443
rect 2141 424 2147 436
rect 1757 277 1779 283
rect 1620 257 1667 263
rect 1645 237 1715 243
rect 1165 144 1171 176
rect 1245 144 1251 196
rect 1277 144 1283 196
rect 1293 164 1299 196
rect 1357 184 1363 236
rect 1373 163 1379 236
rect 1373 157 1388 163
rect 1133 104 1139 136
rect 1229 104 1235 136
rect 1245 124 1251 136
rect 1293 124 1299 136
rect 1277 104 1283 116
rect 1325 104 1331 136
rect 1373 124 1379 136
rect 845 97 899 103
rect 1021 84 1027 96
rect 1165 83 1171 96
rect 1357 84 1363 116
rect 1389 104 1395 156
rect 1485 144 1491 156
rect 1501 124 1507 136
rect 1517 124 1523 196
rect 1549 184 1555 236
rect 1565 124 1571 156
rect 1645 144 1651 237
rect 1709 224 1715 237
rect 1661 143 1667 216
rect 1693 144 1699 216
rect 1709 164 1715 176
rect 1661 137 1683 143
rect 1405 104 1411 116
rect 1453 104 1459 116
rect 1453 84 1459 96
rect 1581 84 1587 116
rect 1140 77 1171 83
rect 1613 43 1619 136
rect 1677 123 1683 137
rect 1725 143 1731 176
rect 1757 164 1763 277
rect 1981 277 2019 283
rect 1789 164 1795 276
rect 1885 263 1891 276
rect 1933 263 1939 276
rect 1981 263 1987 277
rect 1885 257 1939 263
rect 1965 257 1987 263
rect 1965 243 1971 257
rect 2013 244 2019 277
rect 2029 264 2035 296
rect 2061 264 2067 276
rect 2141 264 2147 416
rect 2237 344 2243 416
rect 2189 304 2195 336
rect 2237 304 2243 316
rect 2189 284 2195 296
rect 2253 284 2259 416
rect 2269 284 2275 437
rect 2317 424 2323 436
rect 2333 403 2339 456
rect 2461 444 2467 537
rect 2493 524 2499 536
rect 2493 504 2499 516
rect 2317 397 2339 403
rect 2317 384 2323 397
rect 2333 323 2339 336
rect 2333 317 2355 323
rect 2349 303 2355 317
rect 2397 304 2403 396
rect 2493 324 2499 496
rect 2349 297 2364 303
rect 2509 284 2515 557
rect 2525 524 2531 536
rect 2397 277 2428 283
rect 1917 237 1971 243
rect 1917 224 1923 237
rect 1981 224 1987 236
rect 1892 217 1907 223
rect 1901 203 1907 217
rect 2029 217 2067 223
rect 1933 203 1939 216
rect 1901 197 1939 203
rect 1837 164 1843 196
rect 1709 137 1731 143
rect 1709 123 1715 137
rect 1677 117 1715 123
rect 1549 37 1619 43
rect 1549 24 1555 37
rect 1645 24 1651 116
rect 1901 103 1907 116
rect 1949 104 1955 116
rect 1885 97 1907 103
rect 1885 84 1891 97
rect 1933 84 1939 96
rect 1965 83 1971 216
rect 1981 164 1987 176
rect 1981 104 1987 156
rect 2029 124 2035 217
rect 2045 164 2051 196
rect 2061 184 2067 217
rect 2061 104 2067 156
rect 2077 124 2083 256
rect 2157 204 2163 236
rect 2173 183 2179 196
rect 2093 177 2179 183
rect 2093 164 2099 177
rect 2253 164 2259 236
rect 2125 157 2163 163
rect 2125 143 2131 157
rect 2157 144 2163 157
rect 2221 144 2227 156
rect 2109 137 2131 143
rect 2004 97 2051 103
rect 1965 77 2019 83
rect 2013 63 2019 77
rect 2045 83 2051 97
rect 2093 84 2099 96
rect 2045 77 2083 83
rect 2077 63 2083 77
rect 2109 63 2115 137
rect 2141 124 2147 136
rect 2253 124 2259 156
rect 2269 143 2275 256
rect 2397 224 2403 277
rect 2525 264 2531 436
rect 2541 344 2547 636
rect 2557 624 2563 656
rect 2589 624 2595 677
rect 2573 524 2579 616
rect 2589 524 2595 596
rect 2605 584 2611 736
rect 2621 564 2627 596
rect 2621 544 2627 556
rect 2637 544 2643 877
rect 2669 704 2675 996
rect 2685 903 2691 1057
rect 2701 924 2707 1117
rect 2765 1103 2771 1316
rect 2733 1097 2771 1103
rect 2733 1084 2739 1097
rect 2733 924 2739 1036
rect 2749 984 2755 1076
rect 2765 1044 2771 1076
rect 2685 897 2707 903
rect 2701 863 2707 897
rect 2724 897 2739 903
rect 2685 857 2707 863
rect 2733 863 2739 897
rect 2733 857 2755 863
rect 2685 704 2691 857
rect 2749 803 2755 857
rect 2781 823 2787 1276
rect 2797 1204 2803 1316
rect 2813 1284 2819 1316
rect 2797 1044 2803 1096
rect 2813 964 2819 1196
rect 2829 1084 2835 1136
rect 2861 1083 2867 1276
rect 2852 1077 2867 1083
rect 2836 1057 2860 1063
rect 2829 957 2844 963
rect 2804 837 2819 843
rect 2781 817 2803 823
rect 2749 797 2780 803
rect 2717 724 2723 776
rect 2701 684 2707 696
rect 2653 564 2659 676
rect 2701 584 2707 616
rect 2749 544 2755 797
rect 2765 704 2771 756
rect 2781 684 2787 716
rect 2765 664 2771 676
rect 2797 663 2803 817
rect 2813 804 2819 837
rect 2829 744 2835 957
rect 2877 944 2883 1096
rect 2893 1044 2899 1436
rect 2909 1384 2915 1637
rect 2925 1604 2931 1616
rect 2925 1524 2931 1596
rect 3181 1584 3187 1856
rect 3197 1784 3203 1877
rect 3213 1864 3219 1876
rect 3229 1843 3235 2117
rect 3245 2084 3251 2536
rect 3277 2063 3283 2597
rect 3309 2544 3315 2576
rect 3325 2564 3331 2636
rect 3357 2584 3363 2656
rect 3405 2604 3411 2696
rect 3453 2684 3459 2716
rect 3469 2664 3475 2757
rect 3517 2737 3555 2743
rect 3517 2724 3523 2737
rect 3549 2724 3555 2737
rect 3533 2684 3539 2716
rect 3453 2564 3459 2616
rect 3485 2604 3491 2676
rect 3501 2624 3507 2656
rect 3517 2624 3523 2636
rect 3325 2404 3331 2536
rect 3293 2304 3299 2376
rect 3341 2344 3347 2536
rect 3373 2464 3379 2536
rect 3453 2444 3459 2516
rect 3469 2484 3475 2596
rect 3485 2484 3491 2576
rect 3501 2544 3507 2576
rect 3485 2463 3491 2476
rect 3469 2457 3491 2463
rect 3389 2384 3395 2436
rect 3325 2317 3379 2323
rect 3325 2304 3331 2317
rect 3373 2304 3379 2317
rect 3309 2244 3315 2256
rect 3341 2244 3347 2276
rect 3357 2104 3363 2296
rect 3373 2224 3379 2276
rect 3389 2184 3395 2336
rect 3421 2284 3427 2436
rect 3469 2423 3475 2457
rect 3533 2444 3539 2636
rect 3565 2604 3571 2756
rect 3597 2684 3603 2716
rect 3613 2684 3619 2836
rect 3661 2784 3667 2836
rect 3693 2723 3699 2836
rect 3773 2804 3779 3056
rect 3805 2983 3811 3056
rect 3837 3044 3843 3057
rect 3869 3044 3875 3057
rect 3901 2984 3907 3077
rect 3789 2977 3811 2983
rect 3789 2924 3795 2977
rect 3805 2864 3811 2936
rect 3828 2917 3859 2923
rect 3853 2904 3859 2917
rect 3837 2804 3843 2836
rect 3853 2804 3859 2896
rect 3869 2864 3875 2956
rect 3901 2903 3907 2916
rect 3917 2904 3923 2936
rect 3965 2924 3971 2936
rect 4020 2917 4028 2923
rect 3949 2904 3955 2916
rect 3885 2897 3907 2903
rect 3885 2804 3891 2897
rect 3901 2784 3907 2796
rect 3693 2717 3731 2723
rect 3725 2704 3731 2717
rect 3677 2664 3683 2676
rect 3693 2664 3699 2696
rect 3741 2683 3747 2756
rect 3757 2704 3763 2756
rect 3773 2684 3779 2776
rect 3789 2704 3795 2716
rect 4013 2704 4019 2876
rect 4045 2784 4051 3096
rect 4077 2984 4083 3076
rect 4093 2984 4099 3097
rect 4109 2956 4115 3036
rect 4061 2883 4067 2936
rect 4093 2884 4099 2916
rect 4061 2877 4083 2883
rect 3725 2677 3747 2683
rect 3565 2503 3571 2576
rect 3613 2544 3619 2636
rect 3725 2604 3731 2677
rect 3565 2497 3587 2503
rect 3581 2444 3587 2497
rect 3453 2417 3475 2423
rect 3453 2244 3459 2417
rect 3517 2397 3587 2403
rect 3517 2288 3523 2397
rect 3581 2383 3587 2397
rect 3581 2377 3612 2383
rect 3629 2343 3635 2436
rect 3645 2364 3651 2536
rect 3661 2523 3667 2596
rect 3757 2584 3763 2656
rect 3805 2604 3811 2676
rect 3821 2604 3827 2696
rect 3661 2517 3683 2523
rect 3677 2444 3683 2517
rect 3693 2504 3699 2556
rect 3789 2484 3795 2536
rect 3837 2504 3843 2556
rect 3853 2544 3859 2596
rect 3885 2584 3891 2656
rect 3917 2524 3923 2656
rect 3997 2584 4003 2616
rect 4013 2564 4019 2656
rect 3933 2544 3939 2556
rect 3661 2424 3667 2436
rect 3661 2403 3667 2416
rect 3661 2397 3683 2403
rect 3581 2337 3635 2343
rect 3549 2264 3555 2276
rect 3373 2124 3379 2156
rect 3421 2144 3427 2236
rect 3469 2144 3475 2216
rect 3517 2184 3523 2236
rect 3565 2184 3571 2296
rect 3581 2143 3587 2337
rect 3597 2264 3603 2316
rect 3677 2304 3683 2397
rect 3741 2284 3747 2416
rect 3693 2264 3699 2276
rect 3661 2244 3667 2256
rect 3725 2244 3731 2256
rect 3757 2243 3763 2476
rect 3853 2444 3859 2516
rect 3869 2464 3875 2516
rect 3885 2484 3891 2496
rect 3933 2483 3939 2536
rect 3917 2477 3939 2483
rect 3837 2384 3843 2436
rect 3917 2404 3923 2477
rect 3981 2444 3987 2476
rect 3940 2437 3964 2443
rect 3997 2404 4003 2556
rect 4029 2444 4035 2676
rect 4045 2544 4051 2696
rect 4061 2564 4067 2856
rect 4077 2803 4083 2877
rect 4077 2797 4099 2803
rect 4045 2423 4051 2516
rect 4029 2417 4051 2423
rect 4029 2404 4035 2417
rect 3828 2337 3891 2343
rect 3869 2304 3875 2316
rect 3821 2264 3827 2296
rect 3885 2284 3891 2337
rect 3853 2264 3859 2276
rect 3901 2264 3907 2376
rect 3917 2304 3923 2336
rect 4061 2304 4067 2516
rect 4077 2504 4083 2736
rect 4093 2524 4099 2797
rect 4125 2683 4131 2916
rect 4157 2804 4163 3116
rect 4205 3024 4211 3096
rect 4285 3024 4291 3056
rect 4292 3017 4307 3023
rect 4285 2944 4291 2976
rect 4237 2743 4243 2776
rect 4237 2737 4259 2743
rect 4109 2677 4131 2683
rect 4109 2664 4115 2677
rect 4141 2544 4147 2676
rect 4173 2584 4179 2636
rect 4237 2624 4243 2676
rect 4237 2604 4243 2616
rect 4109 2537 4124 2543
rect 4109 2524 4115 2537
rect 4205 2524 4211 2576
rect 4253 2524 4259 2737
rect 4269 2543 4275 2676
rect 4285 2564 4291 2756
rect 4269 2537 4291 2543
rect 3997 2302 4003 2303
rect 3997 2284 4003 2294
rect 3757 2237 3779 2243
rect 3693 2184 3699 2216
rect 3565 2137 3587 2143
rect 3501 2124 3507 2136
rect 3533 2124 3539 2136
rect 3565 2124 3571 2137
rect 3629 2124 3635 2136
rect 3645 2124 3651 2156
rect 3588 2117 3603 2123
rect 3245 2057 3283 2063
rect 3245 1924 3251 2057
rect 3261 2024 3267 2036
rect 3261 1884 3267 1936
rect 3277 1924 3283 1996
rect 3277 1884 3283 1916
rect 3293 1884 3299 2016
rect 3325 1924 3331 2096
rect 3341 1924 3347 1976
rect 3357 1944 3363 2056
rect 3229 1837 3267 1843
rect 3213 1764 3219 1836
rect 3261 1824 3267 1837
rect 3229 1684 3235 1716
rect 3245 1703 3251 1816
rect 3277 1784 3283 1856
rect 3293 1804 3299 1816
rect 3293 1724 3299 1796
rect 3309 1744 3315 1836
rect 3325 1824 3331 1916
rect 3357 1843 3363 1896
rect 3373 1864 3379 1996
rect 3453 1984 3459 2116
rect 3549 2004 3555 2036
rect 3597 2004 3603 2117
rect 3709 2103 3715 2236
rect 3700 2097 3715 2103
rect 3405 1884 3411 1896
rect 3389 1863 3395 1876
rect 3389 1857 3404 1863
rect 3357 1837 3395 1843
rect 3389 1823 3395 1837
rect 3389 1817 3411 1823
rect 3325 1784 3331 1796
rect 3357 1764 3363 1796
rect 3373 1764 3379 1816
rect 3389 1784 3395 1796
rect 3405 1764 3411 1817
rect 3421 1804 3427 1936
rect 3581 1924 3587 1996
rect 3613 1964 3619 2096
rect 3645 2017 3683 2023
rect 3533 1903 3539 1916
rect 3524 1897 3539 1903
rect 3437 1884 3443 1896
rect 3549 1884 3555 1896
rect 3565 1884 3571 1896
rect 3597 1864 3603 1896
rect 3437 1804 3443 1856
rect 3389 1724 3395 1756
rect 3245 1697 3315 1703
rect 3245 1677 3260 1683
rect 3213 1663 3219 1676
rect 3245 1663 3251 1677
rect 3213 1657 3251 1663
rect 3277 1563 3283 1676
rect 3245 1557 3283 1563
rect 3245 1544 3251 1557
rect 2957 1537 2988 1543
rect 2957 1523 2963 1537
rect 2941 1517 2963 1523
rect 2941 1504 2947 1517
rect 3021 1503 3027 1516
rect 3101 1504 3107 1536
rect 3117 1504 3123 1536
rect 3140 1517 3171 1523
rect 3021 1497 3059 1503
rect 2941 1464 2947 1476
rect 3005 1464 3011 1496
rect 2925 1283 2931 1336
rect 2909 1277 2931 1283
rect 2845 864 2851 916
rect 2861 904 2867 936
rect 2893 924 2899 1036
rect 2909 944 2915 1277
rect 2941 1224 2947 1436
rect 2989 1384 2995 1456
rect 2989 1344 2995 1356
rect 3005 1324 3011 1416
rect 3053 1364 3059 1497
rect 3165 1503 3171 1517
rect 3236 1517 3251 1523
rect 3156 1497 3171 1503
rect 3172 1457 3187 1463
rect 3101 1444 3107 1456
rect 3069 1343 3075 1396
rect 3085 1364 3091 1436
rect 3112 1406 3113 1414
rect 3121 1406 3123 1414
rect 3131 1406 3133 1414
rect 3141 1406 3143 1414
rect 3151 1406 3160 1414
rect 3181 1404 3187 1457
rect 3197 1444 3203 1476
rect 3245 1384 3251 1517
rect 3261 1504 3267 1536
rect 3277 1484 3283 1557
rect 3309 1484 3315 1697
rect 3341 1502 3347 1503
rect 3117 1343 3123 1356
rect 3069 1337 3123 1343
rect 2973 1304 2979 1316
rect 3021 1263 3027 1276
rect 3021 1257 3107 1263
rect 2925 1044 2931 1096
rect 2925 904 2931 916
rect 2925 864 2931 896
rect 2941 864 2947 1116
rect 2973 1104 2979 1216
rect 3053 1144 3059 1236
rect 3021 1104 3027 1136
rect 2957 944 2963 1056
rect 2973 1024 2979 1096
rect 3069 1084 3075 1156
rect 3085 1144 3091 1176
rect 3101 1103 3107 1257
rect 3117 1124 3123 1236
rect 3133 1184 3139 1376
rect 3149 1204 3155 1376
rect 3165 1284 3171 1336
rect 3245 1324 3251 1336
rect 3181 1304 3187 1316
rect 3165 1104 3171 1196
rect 3181 1184 3187 1276
rect 3213 1204 3219 1236
rect 3101 1097 3116 1103
rect 3085 1084 3091 1096
rect 3101 1063 3107 1076
rect 3085 1057 3107 1063
rect 2973 924 2979 956
rect 3005 944 3011 1036
rect 3021 984 3027 1016
rect 2989 924 2995 936
rect 2989 863 2995 896
rect 3021 884 3027 916
rect 3037 883 3043 976
rect 3053 944 3059 1056
rect 3069 964 3075 1036
rect 3085 1024 3091 1057
rect 3172 1037 3187 1043
rect 3112 1006 3113 1014
rect 3121 1006 3123 1014
rect 3131 1006 3133 1014
rect 3141 1006 3143 1014
rect 3151 1006 3160 1014
rect 3085 944 3091 996
rect 3101 923 3107 956
rect 3092 917 3107 923
rect 3069 904 3075 916
rect 3037 877 3059 883
rect 3005 863 3011 876
rect 3053 864 3059 877
rect 3085 864 3091 876
rect 2989 857 3011 863
rect 2909 843 2915 856
rect 2941 843 2947 856
rect 2909 837 2947 843
rect 2845 784 2851 796
rect 2813 664 2819 676
rect 2781 657 2803 663
rect 2781 644 2787 657
rect 2829 544 2835 716
rect 2925 704 2931 716
rect 2941 704 2947 816
rect 2973 723 2979 856
rect 3101 844 3107 876
rect 3117 823 3123 836
rect 3069 817 3123 823
rect 3069 804 3075 817
rect 3021 763 3027 796
rect 3085 783 3091 796
rect 3053 777 3091 783
rect 3053 763 3059 777
rect 3021 757 3059 763
rect 2973 717 2995 723
rect 2989 704 2995 717
rect 2845 697 2860 703
rect 2845 584 2851 697
rect 2861 624 2867 656
rect 2877 604 2883 676
rect 2973 664 2979 696
rect 2973 644 2979 656
rect 2621 483 2627 516
rect 2637 504 2643 516
rect 2781 504 2787 536
rect 2893 524 2899 616
rect 2973 543 2979 636
rect 2964 537 2979 543
rect 2909 524 2915 536
rect 2653 483 2659 496
rect 2813 484 2819 496
rect 2621 477 2659 483
rect 2829 463 2835 516
rect 2813 457 2835 463
rect 2733 437 2748 443
rect 2557 304 2563 436
rect 2573 283 2579 336
rect 2605 324 2611 436
rect 2621 357 2691 363
rect 2621 344 2627 357
rect 2557 277 2579 283
rect 2413 224 2419 236
rect 2413 184 2419 216
rect 2429 184 2435 256
rect 2541 184 2547 236
rect 2557 224 2563 277
rect 2596 257 2620 263
rect 2573 224 2579 236
rect 2653 223 2659 276
rect 2669 264 2675 316
rect 2685 224 2691 357
rect 2717 304 2723 356
rect 2733 344 2739 437
rect 2813 423 2819 457
rect 2756 417 2819 423
rect 2829 344 2835 436
rect 2893 403 2899 516
rect 2909 504 2915 516
rect 2989 463 2995 536
rect 3005 524 3011 736
rect 3037 703 3043 716
rect 3021 697 3043 703
rect 3021 624 3027 697
rect 3069 564 3075 676
rect 3085 664 3091 736
rect 3133 724 3139 956
rect 3101 664 3107 696
rect 3133 684 3139 716
rect 3181 704 3187 1037
rect 3197 924 3203 1176
rect 3261 1124 3267 1476
rect 3277 1344 3283 1476
rect 3341 1464 3347 1494
rect 3373 1404 3379 1716
rect 3437 1544 3443 1736
rect 3453 1484 3459 1576
rect 3469 1564 3475 1816
rect 3565 1744 3571 1756
rect 3508 1737 3523 1743
rect 3501 1663 3507 1716
rect 3485 1657 3507 1663
rect 3300 1397 3331 1403
rect 3325 1384 3331 1397
rect 3389 1363 3395 1416
rect 3453 1404 3459 1456
rect 3389 1357 3411 1363
rect 3277 1324 3283 1336
rect 3293 1324 3299 1336
rect 3293 1144 3299 1256
rect 3293 1084 3299 1096
rect 3309 1084 3315 1136
rect 3245 1004 3251 1076
rect 3293 944 3299 1056
rect 3341 944 3347 1296
rect 3405 1283 3411 1357
rect 3421 1304 3427 1376
rect 3405 1277 3427 1283
rect 3373 1104 3379 1276
rect 3373 1084 3379 1096
rect 3389 984 3395 1256
rect 3405 1024 3411 1116
rect 3421 1103 3427 1277
rect 3437 1123 3443 1396
rect 3485 1284 3491 1657
rect 3517 1444 3523 1737
rect 3533 1604 3539 1736
rect 3581 1724 3587 1776
rect 3597 1723 3603 1836
rect 3613 1764 3619 1876
rect 3629 1843 3635 2016
rect 3645 1924 3651 2017
rect 3677 2004 3683 2017
rect 3661 1983 3667 1996
rect 3661 1977 3692 1983
rect 3741 1983 3747 2236
rect 3757 2164 3763 2216
rect 3757 2144 3763 2156
rect 3773 2104 3779 2237
rect 3789 2124 3795 2136
rect 3805 2103 3811 2116
rect 3789 2097 3811 2103
rect 3789 1984 3795 2097
rect 3709 1977 3747 1983
rect 3709 1944 3715 1977
rect 3725 1957 3779 1963
rect 3725 1944 3731 1957
rect 3677 1904 3683 1936
rect 3741 1924 3747 1936
rect 3725 1864 3731 1896
rect 3757 1883 3763 1916
rect 3773 1904 3779 1957
rect 3757 1877 3779 1883
rect 3629 1837 3651 1843
rect 3613 1743 3619 1756
rect 3613 1737 3628 1743
rect 3645 1724 3651 1837
rect 3661 1804 3667 1856
rect 3597 1717 3619 1723
rect 3565 1584 3571 1716
rect 3613 1704 3619 1717
rect 3581 1604 3587 1636
rect 3549 1563 3555 1576
rect 3549 1557 3571 1563
rect 3565 1504 3571 1557
rect 3613 1504 3619 1596
rect 3629 1504 3635 1596
rect 3629 1464 3635 1476
rect 3437 1117 3459 1123
rect 3453 1104 3459 1117
rect 3501 1104 3507 1316
rect 3421 1097 3443 1103
rect 3373 964 3379 976
rect 3213 924 3219 936
rect 3389 924 3395 956
rect 3245 844 3251 916
rect 3213 803 3219 836
rect 3197 797 3219 803
rect 3197 704 3203 797
rect 3309 744 3315 916
rect 3149 643 3155 656
rect 3149 637 3187 643
rect 3085 543 3091 636
rect 3112 606 3113 614
rect 3121 606 3123 614
rect 3131 606 3133 614
rect 3141 606 3143 614
rect 3151 606 3160 614
rect 3181 604 3187 637
rect 3117 564 3123 576
rect 3085 537 3100 543
rect 3021 524 3027 536
rect 3012 497 3036 503
rect 3117 463 3123 516
rect 2989 457 3011 463
rect 3005 443 3011 457
rect 3053 457 3123 463
rect 3053 443 3059 457
rect 3005 437 3059 443
rect 2973 404 2979 436
rect 2893 397 2908 403
rect 2909 377 2995 383
rect 2772 337 2796 343
rect 2717 284 2723 296
rect 2733 284 2739 336
rect 2813 323 2819 336
rect 2797 317 2819 323
rect 2765 304 2771 316
rect 2749 283 2755 296
rect 2797 283 2803 317
rect 2749 277 2803 283
rect 2813 297 2844 303
rect 2701 263 2707 276
rect 2701 257 2732 263
rect 2813 263 2819 297
rect 2877 264 2883 336
rect 2909 304 2915 377
rect 2941 357 2979 363
rect 2941 344 2947 357
rect 2973 344 2979 357
rect 2989 343 2995 377
rect 2989 337 3011 343
rect 2957 324 2963 336
rect 3005 323 3011 337
rect 3037 337 3091 343
rect 3005 317 3027 323
rect 2925 304 2931 316
rect 2989 297 3004 303
rect 2973 284 2979 296
rect 2804 257 2819 263
rect 2909 263 2915 276
rect 2989 263 2995 297
rect 3021 284 3027 317
rect 3037 263 3043 337
rect 3069 284 3075 316
rect 3085 284 3091 337
rect 3133 324 3139 556
rect 3165 544 3171 576
rect 3197 543 3203 696
rect 3213 684 3219 696
rect 3229 644 3235 676
rect 3245 663 3251 716
rect 3293 663 3299 696
rect 3245 657 3267 663
rect 3229 584 3235 616
rect 3245 564 3251 636
rect 3261 624 3267 657
rect 3277 657 3299 663
rect 3188 537 3203 543
rect 3181 517 3196 523
rect 3181 504 3187 517
rect 3149 404 3155 496
rect 3229 464 3235 556
rect 3277 543 3283 657
rect 3293 564 3299 636
rect 3309 543 3315 716
rect 3325 644 3331 696
rect 3341 684 3347 896
rect 3405 884 3411 1016
rect 3405 724 3411 876
rect 3421 764 3427 976
rect 3437 884 3443 1097
rect 3517 1084 3523 1116
rect 3533 1104 3539 1276
rect 3565 1224 3571 1436
rect 3629 1364 3635 1376
rect 3597 1283 3603 1316
rect 3581 1277 3603 1283
rect 3469 1024 3475 1076
rect 3565 1064 3571 1196
rect 3581 1184 3587 1277
rect 3581 1104 3587 1176
rect 3485 1024 3491 1036
rect 3517 1004 3523 1056
rect 3549 1044 3555 1056
rect 3501 964 3507 976
rect 3565 964 3571 1056
rect 3597 1044 3603 1056
rect 3661 1044 3667 1796
rect 3741 1783 3747 1856
rect 3757 1784 3763 1796
rect 3725 1777 3747 1783
rect 3677 1364 3683 1756
rect 3693 1744 3699 1756
rect 3693 1504 3699 1716
rect 3725 1704 3731 1777
rect 3773 1764 3779 1877
rect 3789 1863 3795 1916
rect 3805 1904 3811 1996
rect 3837 1984 3843 2156
rect 3853 2124 3859 2136
rect 3869 2124 3875 2136
rect 3885 2124 3891 2196
rect 3821 1923 3827 1976
rect 3853 1944 3859 2116
rect 3821 1917 3859 1923
rect 3853 1903 3859 1917
rect 3885 1923 3891 2116
rect 3876 1917 3891 1923
rect 3853 1897 3868 1903
rect 3789 1857 3827 1863
rect 3741 1724 3747 1756
rect 3821 1743 3827 1857
rect 3837 1804 3843 1896
rect 3901 1824 3907 2176
rect 3917 2124 3923 2156
rect 3924 2097 3932 2103
rect 3949 2063 3955 2136
rect 3965 2104 3971 2116
rect 3981 2104 3987 2116
rect 4061 2104 4067 2118
rect 3997 2064 4003 2096
rect 3933 2057 3955 2063
rect 3933 1923 3939 2057
rect 3956 1977 3964 1983
rect 3933 1917 3964 1923
rect 3933 1904 3939 1917
rect 3981 1904 3987 1916
rect 3997 1884 4003 1976
rect 4013 1884 4019 2056
rect 4029 1984 4035 2036
rect 4045 1964 4051 1996
rect 4045 1924 4051 1956
rect 4045 1904 4051 1916
rect 4061 1884 4067 1956
rect 3853 1743 3859 1796
rect 3901 1744 3907 1756
rect 3933 1744 3939 1876
rect 4013 1857 4028 1863
rect 4013 1764 4019 1857
rect 3805 1737 3843 1743
rect 3853 1737 3875 1743
rect 3725 1564 3731 1696
rect 3709 1537 3724 1543
rect 3709 1504 3715 1537
rect 3757 1384 3763 1636
rect 3805 1444 3811 1737
rect 3837 1724 3843 1737
rect 3869 1723 3875 1737
rect 3869 1717 3884 1723
rect 3821 1703 3827 1716
rect 3965 1704 3971 1718
rect 3821 1697 3852 1703
rect 3933 1683 3939 1696
rect 3981 1683 3987 1756
rect 3917 1677 3939 1683
rect 3965 1677 3987 1683
rect 3917 1663 3923 1677
rect 3892 1657 3923 1663
rect 3965 1583 3971 1677
rect 4013 1624 4019 1676
rect 3901 1577 3971 1583
rect 3901 1564 3907 1577
rect 3949 1557 3987 1563
rect 3949 1543 3955 1557
rect 3933 1537 3955 1543
rect 3933 1524 3939 1537
rect 3981 1524 3987 1557
rect 3949 1504 3955 1516
rect 3853 1502 3859 1503
rect 3853 1484 3859 1494
rect 3917 1484 3923 1496
rect 4013 1484 4019 1496
rect 4029 1484 4035 1836
rect 4045 1824 4051 1876
rect 4045 1584 4051 1616
rect 4077 1503 4083 2096
rect 4093 1964 4099 2436
rect 4125 2384 4131 2516
rect 4253 2504 4259 2516
rect 4269 2444 4275 2516
rect 4285 2504 4291 2537
rect 4301 2524 4307 3017
rect 4317 2984 4323 3056
rect 4397 3044 4403 3117
rect 4429 3104 4435 3116
rect 4413 3064 4419 3076
rect 4461 3044 4467 3076
rect 4477 3064 4483 3256
rect 4509 3184 4515 3196
rect 4525 3104 4531 3136
rect 4525 3064 4531 3096
rect 4317 2904 4323 2936
rect 4349 2924 4355 3016
rect 4381 2964 4387 3036
rect 4493 3024 4499 3036
rect 4509 2984 4515 3036
rect 4125 2324 4131 2336
rect 4189 2324 4195 2336
rect 4157 2284 4163 2296
rect 4237 2284 4243 2436
rect 4285 2424 4291 2496
rect 4301 2424 4307 2436
rect 4317 2403 4323 2656
rect 4349 2544 4355 2696
rect 4381 2684 4387 2936
rect 4525 2924 4531 2936
rect 4557 2904 4563 2936
rect 4573 2924 4579 2956
rect 4605 2903 4611 2956
rect 4637 2944 4643 3276
rect 4664 3206 4665 3214
rect 4673 3206 4675 3214
rect 4683 3206 4685 3214
rect 4693 3206 4695 3214
rect 4703 3206 4712 3214
rect 4669 3102 4675 3136
rect 4733 3084 4739 3336
rect 4765 3084 4771 3357
rect 4797 3324 4803 3496
rect 4861 3483 4867 3496
rect 4852 3477 4867 3483
rect 4852 3337 4867 3343
rect 4861 3324 4867 3337
rect 4781 3124 4787 3316
rect 4845 3304 4851 3316
rect 4893 3184 4899 3296
rect 4781 3104 4787 3116
rect 4877 3084 4883 3096
rect 4605 2897 4620 2903
rect 4605 2743 4611 2897
rect 4653 2884 4659 2956
rect 4733 2944 4739 3036
rect 4685 2844 4691 2936
rect 4733 2924 4739 2936
rect 4893 2884 4899 3036
rect 4909 2944 4915 3716
rect 5149 3704 5155 3716
rect 5165 3644 5171 3756
rect 5245 3744 5251 3756
rect 4964 3497 4972 3503
rect 5085 3484 5091 3636
rect 5181 3524 5187 3636
rect 5197 3584 5203 3696
rect 5229 3584 5235 3616
rect 5245 3544 5251 3736
rect 5277 3723 5283 3796
rect 5277 3717 5292 3723
rect 5309 3604 5315 3836
rect 5357 3724 5363 3836
rect 5373 3764 5379 3856
rect 5373 3724 5379 3736
rect 5373 3704 5379 3716
rect 5325 3624 5331 3696
rect 5357 3683 5363 3696
rect 5389 3683 5395 3716
rect 5357 3677 5395 3683
rect 5357 3584 5363 3616
rect 5421 3584 5427 3816
rect 5453 3804 5459 3856
rect 5517 3764 5523 3836
rect 5677 3784 5683 3816
rect 5725 3803 5731 3876
rect 5725 3797 5740 3803
rect 5741 3784 5747 3796
rect 5661 3764 5667 3776
rect 5437 3704 5443 3716
rect 5117 3504 5123 3516
rect 5021 3364 5027 3456
rect 5117 3424 5123 3436
rect 5197 3384 5203 3516
rect 5229 3404 5235 3496
rect 5261 3484 5267 3496
rect 5277 3484 5283 3576
rect 5277 3464 5283 3476
rect 5277 3384 5283 3436
rect 5293 3404 5299 3436
rect 4957 3324 4963 3336
rect 5021 3084 5027 3356
rect 5245 3344 5251 3356
rect 5293 3344 5299 3356
rect 5053 3104 5059 3316
rect 5085 3304 5091 3336
rect 5117 3324 5123 3336
rect 5245 3304 5251 3336
rect 5309 3324 5315 3536
rect 5325 3504 5331 3576
rect 5373 3524 5379 3536
rect 5421 3504 5427 3576
rect 5469 3504 5475 3676
rect 5485 3664 5491 3756
rect 5757 3744 5763 4016
rect 5789 4004 5795 4136
rect 5789 3964 5795 3996
rect 5837 3924 5843 4116
rect 5853 4104 5859 4196
rect 5901 4124 5907 4276
rect 5917 4244 5923 4296
rect 5933 4284 5939 4296
rect 5949 4264 5955 4296
rect 5988 4277 6003 4283
rect 5981 4244 5987 4256
rect 5997 4224 6003 4277
rect 6013 4203 6019 4256
rect 6029 4204 6035 4356
rect 5997 4197 6019 4203
rect 5917 4144 5923 4196
rect 5949 4184 5955 4196
rect 5853 4024 5859 4096
rect 5885 4004 5891 4116
rect 5917 4104 5923 4116
rect 5933 4084 5939 4136
rect 5981 4124 5987 4156
rect 5997 4104 6003 4197
rect 6061 4184 6067 4276
rect 6077 4184 6083 4376
rect 6093 4264 6099 4276
rect 6109 4163 6115 4477
rect 6125 4344 6131 4436
rect 6141 4323 6147 4436
rect 6157 4384 6163 4416
rect 6173 4364 6179 4496
rect 6189 4444 6195 4536
rect 6205 4504 6211 4516
rect 6237 4424 6243 4496
rect 6285 4464 6291 4536
rect 6132 4317 6147 4323
rect 6093 4157 6115 4163
rect 6061 4144 6067 4156
rect 5853 3984 5859 3996
rect 5901 3984 5907 4036
rect 5949 3984 5955 4016
rect 5885 3904 5891 3936
rect 5773 3884 5779 3896
rect 5789 3884 5795 3896
rect 5869 3884 5875 3896
rect 5901 3883 5907 3936
rect 5933 3884 5939 3956
rect 5885 3877 5907 3883
rect 5789 3844 5795 3876
rect 5869 3864 5875 3876
rect 5853 3823 5859 3836
rect 5853 3817 5875 3823
rect 5517 3737 5532 3743
rect 5517 3724 5523 3737
rect 5629 3724 5635 3736
rect 5725 3724 5731 3736
rect 5757 3704 5763 3716
rect 5684 3697 5724 3703
rect 5517 3644 5523 3696
rect 5549 3664 5555 3676
rect 5581 3643 5587 3696
rect 5677 3684 5683 3696
rect 5773 3664 5779 3736
rect 5565 3637 5603 3643
rect 5501 3624 5507 3636
rect 5565 3624 5571 3637
rect 5597 3624 5603 3637
rect 5581 3584 5587 3616
rect 5469 3484 5475 3496
rect 5485 3484 5491 3496
rect 5549 3484 5555 3556
rect 5645 3523 5651 3636
rect 5757 3584 5763 3656
rect 5645 3517 5699 3523
rect 5565 3504 5571 3516
rect 5629 3504 5635 3516
rect 5693 3504 5699 3517
rect 5581 3483 5587 3496
rect 5661 3484 5667 3496
rect 5677 3484 5683 3496
rect 5572 3477 5587 3483
rect 5693 3477 5724 3483
rect 5325 3424 5331 3476
rect 5421 3444 5427 3476
rect 5453 3404 5459 3436
rect 5389 3344 5395 3356
rect 5437 3344 5443 3376
rect 5325 3337 5363 3343
rect 5325 3324 5331 3337
rect 5341 3304 5347 3316
rect 5357 3304 5363 3337
rect 5444 3337 5459 3343
rect 5421 3324 5427 3336
rect 5380 3317 5395 3323
rect 5389 3244 5395 3317
rect 5453 3323 5459 3337
rect 5453 3317 5484 3323
rect 4973 2964 4979 2976
rect 5021 2924 5027 2936
rect 5021 2884 5027 2896
rect 4621 2764 4627 2836
rect 4605 2737 4627 2743
rect 4397 2704 4403 2736
rect 4477 2684 4483 2696
rect 4445 2664 4451 2676
rect 4333 2524 4339 2536
rect 4333 2444 4339 2516
rect 4301 2397 4323 2403
rect 4276 2377 4284 2383
rect 4141 2264 4147 2276
rect 4253 2264 4259 2376
rect 4285 2264 4291 2276
rect 4253 2184 4259 2256
rect 4109 1924 4115 2056
rect 4125 1924 4131 2156
rect 4269 2144 4275 2156
rect 4237 2064 4243 2136
rect 4253 2104 4259 2116
rect 4285 2104 4291 2236
rect 4301 2144 4307 2397
rect 4349 2324 4355 2336
rect 4365 2284 4371 2516
rect 4397 2504 4403 2656
rect 4493 2604 4499 2696
rect 4429 2524 4435 2596
rect 4477 2564 4483 2596
rect 4509 2583 4515 2616
rect 4493 2577 4515 2583
rect 4445 2444 4451 2536
rect 4461 2524 4467 2536
rect 4477 2503 4483 2516
rect 4461 2497 4483 2503
rect 4381 2284 4387 2296
rect 4356 2277 4364 2283
rect 4333 2084 4339 2096
rect 4157 2004 4163 2056
rect 4189 2023 4195 2036
rect 4189 2017 4211 2023
rect 4125 1917 4128 1924
rect 4093 1824 4099 1916
rect 4157 1884 4163 1996
rect 4173 1917 4188 1923
rect 4173 1904 4179 1917
rect 4205 1903 4211 2017
rect 4221 1937 4252 1943
rect 4221 1924 4227 1937
rect 4269 1923 4275 2036
rect 4301 1944 4307 1956
rect 4253 1917 4275 1923
rect 4205 1897 4227 1903
rect 4125 1784 4131 1856
rect 4100 1777 4115 1783
rect 4109 1744 4115 1777
rect 4109 1623 4115 1676
rect 4141 1624 4147 1816
rect 4205 1744 4211 1876
rect 4221 1784 4227 1897
rect 4237 1884 4243 1916
rect 4253 1904 4259 1917
rect 4237 1804 4243 1876
rect 4269 1724 4275 1896
rect 4285 1724 4291 1796
rect 4189 1704 4195 1716
rect 4240 1696 4243 1703
rect 4109 1617 4131 1623
rect 4125 1524 4131 1617
rect 4164 1517 4179 1523
rect 4068 1497 4083 1503
rect 4173 1503 4179 1517
rect 4173 1497 4195 1503
rect 3940 1477 3948 1483
rect 3677 1244 3683 1316
rect 3693 1304 3699 1316
rect 3725 1224 3731 1296
rect 3789 1144 3795 1336
rect 3725 1084 3731 1136
rect 3821 1104 3827 1236
rect 3837 1083 3843 1156
rect 3828 1077 3843 1083
rect 3613 984 3619 996
rect 3485 943 3491 956
rect 3485 937 3516 943
rect 3549 937 3564 943
rect 3549 924 3555 937
rect 3469 763 3475 896
rect 3501 843 3507 896
rect 3533 863 3539 916
rect 3533 857 3548 863
rect 3565 844 3571 916
rect 3645 864 3651 996
rect 3501 837 3516 843
rect 3437 757 3475 763
rect 3405 704 3411 716
rect 3389 604 3395 696
rect 3437 684 3443 757
rect 3565 743 3571 836
rect 3581 764 3587 836
rect 3565 737 3587 743
rect 3469 684 3475 696
rect 3405 663 3411 676
rect 3405 657 3459 663
rect 3437 603 3443 636
rect 3453 624 3459 657
rect 3501 623 3507 736
rect 3517 704 3523 716
rect 3581 704 3587 737
rect 3597 704 3603 776
rect 3517 684 3523 696
rect 3581 644 3587 696
rect 3613 683 3619 716
rect 3645 704 3651 716
rect 3604 677 3619 683
rect 3661 664 3667 776
rect 3677 724 3683 876
rect 3677 684 3683 716
rect 3492 617 3507 623
rect 3405 597 3443 603
rect 3453 597 3516 603
rect 3373 564 3379 596
rect 3325 557 3340 563
rect 3325 544 3331 557
rect 3245 537 3283 543
rect 3293 537 3315 543
rect 3197 363 3203 456
rect 3197 357 3219 363
rect 3133 284 3139 316
rect 3181 264 3187 356
rect 3197 324 3203 336
rect 3197 284 3203 316
rect 2909 257 2995 263
rect 3021 257 3043 263
rect 2813 224 2819 236
rect 2637 217 2659 223
rect 2445 177 2483 183
rect 2317 144 2323 176
rect 2269 137 2307 143
rect 2125 104 2131 116
rect 2141 104 2147 116
rect 2157 64 2163 76
rect 2205 64 2211 116
rect 2013 57 2067 63
rect 2077 57 2115 63
rect 2061 43 2067 57
rect 2061 37 2131 43
rect 1576 6 1577 14
rect 1585 6 1587 14
rect 1595 6 1597 14
rect 1605 6 1607 14
rect 1615 6 1624 14
rect 1949 -17 1955 22
rect 2125 3 2131 37
rect 2141 24 2147 56
rect 2221 3 2227 116
rect 2269 104 2275 116
rect 2301 83 2307 137
rect 2349 104 2355 176
rect 2445 144 2451 177
rect 2477 163 2483 177
rect 2477 157 2563 163
rect 2557 143 2563 157
rect 2557 137 2579 143
rect 2461 124 2467 136
rect 2253 77 2307 83
rect 2253 43 2259 77
rect 2381 64 2387 116
rect 2477 104 2483 116
rect 2541 104 2547 136
rect 2573 123 2579 137
rect 2573 117 2595 123
rect 2589 104 2595 117
rect 2637 123 2643 217
rect 2765 217 2803 223
rect 2765 204 2771 217
rect 2797 203 2803 217
rect 2797 197 2812 203
rect 2781 164 2787 196
rect 2829 183 2835 216
rect 2893 204 2899 256
rect 2797 177 2835 183
rect 2717 157 2771 163
rect 2660 137 2707 143
rect 2637 117 2691 123
rect 2621 103 2627 116
rect 2621 97 2659 103
rect 2397 84 2403 96
rect 2541 84 2547 96
rect 2125 -3 2227 3
rect 2237 37 2259 43
rect 2237 -17 2243 37
rect 2365 23 2371 56
rect 2573 44 2579 76
rect 2589 37 2620 43
rect 2397 23 2403 36
rect 2365 17 2403 23
rect 2557 23 2563 36
rect 2589 23 2595 37
rect 2557 17 2595 23
rect 2653 23 2659 97
rect 2685 63 2691 117
rect 2701 83 2707 137
rect 2717 104 2723 157
rect 2765 143 2771 157
rect 2797 143 2803 177
rect 2957 144 2963 236
rect 2765 137 2803 143
rect 2733 104 2739 116
rect 2749 104 2755 136
rect 2820 117 2851 123
rect 2813 104 2819 116
rect 2733 84 2739 96
rect 2797 84 2803 96
rect 2829 84 2835 96
rect 2845 84 2851 117
rect 2701 77 2723 83
rect 2717 63 2723 77
rect 2749 63 2755 76
rect 2685 57 2707 63
rect 2717 57 2755 63
rect 2701 43 2707 57
rect 2861 44 2867 136
rect 2909 104 2915 116
rect 3005 84 3011 196
rect 3021 124 3027 257
rect 3037 163 3043 236
rect 3112 206 3113 214
rect 3121 206 3123 214
rect 3131 206 3133 214
rect 3141 206 3143 214
rect 3151 206 3160 214
rect 3085 183 3091 196
rect 3085 177 3123 183
rect 3037 157 3052 163
rect 3037 44 3043 157
rect 3117 144 3123 177
rect 3197 164 3203 216
rect 3213 163 3219 357
rect 3245 344 3251 537
rect 3293 523 3299 537
rect 3373 524 3379 556
rect 3268 517 3299 523
rect 3332 517 3347 523
rect 3261 497 3299 503
rect 3261 464 3267 497
rect 3229 303 3235 336
rect 3277 303 3283 476
rect 3293 363 3299 497
rect 3341 384 3347 517
rect 3405 523 3411 597
rect 3453 563 3459 597
rect 3437 557 3459 563
rect 3389 517 3411 523
rect 3357 504 3363 516
rect 3389 484 3395 517
rect 3421 483 3427 536
rect 3437 524 3443 557
rect 3549 544 3555 636
rect 3565 564 3571 636
rect 3597 544 3603 556
rect 3453 537 3491 543
rect 3453 524 3459 537
rect 3485 504 3491 537
rect 3501 524 3507 536
rect 3613 523 3619 656
rect 3645 564 3651 596
rect 3661 564 3667 576
rect 3629 543 3635 556
rect 3629 537 3651 543
rect 3604 517 3619 523
rect 3421 477 3436 483
rect 3453 464 3459 476
rect 3293 357 3315 363
rect 3229 297 3251 303
rect 3245 283 3251 297
rect 3261 297 3283 303
rect 3261 283 3267 297
rect 3245 277 3267 283
rect 3229 184 3235 196
rect 3245 164 3251 176
rect 3213 157 3235 163
rect 3204 137 3219 143
rect 3053 117 3091 123
rect 3053 104 3059 117
rect 3085 84 3091 117
rect 2701 37 2723 43
rect 2685 23 2691 36
rect 2717 24 2723 37
rect 2653 17 2691 23
rect 2877 23 2883 36
rect 2836 17 2883 23
rect 3181 3 3187 36
rect 3213 24 3219 137
rect 3229 104 3235 157
rect 3261 103 3267 176
rect 3277 144 3283 276
rect 3245 97 3267 103
rect 3245 3 3251 97
rect 3181 -3 3251 3
rect 1949 -23 2243 -17
rect 3245 -37 3251 -17
rect 3293 -37 3299 336
rect 3309 303 3315 357
rect 3325 344 3331 376
rect 3309 297 3331 303
rect 3309 184 3315 276
rect 3325 224 3331 297
rect 3341 284 3347 296
rect 3373 284 3379 436
rect 3485 384 3491 496
rect 3517 484 3523 516
rect 3501 403 3507 436
rect 3501 397 3523 403
rect 3421 304 3427 336
rect 3517 324 3523 397
rect 3613 384 3619 436
rect 3572 337 3580 343
rect 3476 317 3507 323
rect 3341 244 3347 256
rect 3309 164 3315 176
rect 3325 124 3331 156
rect 3341 103 3347 156
rect 3332 97 3347 103
rect 3357 24 3363 236
rect 3421 224 3427 276
rect 3453 123 3459 216
rect 3469 164 3475 296
rect 3485 264 3491 276
rect 3396 117 3443 123
rect 3453 117 3468 123
rect 3437 83 3443 117
rect 3437 77 3475 83
rect 3469 44 3475 77
rect 3501 24 3507 317
rect 3533 303 3539 316
rect 3549 304 3555 336
rect 3645 324 3651 537
rect 3677 483 3683 516
rect 3693 504 3699 976
rect 3709 904 3715 956
rect 3725 944 3731 1076
rect 3805 944 3811 1016
rect 3869 963 3875 1096
rect 3885 1084 3891 1156
rect 3901 1104 3907 1396
rect 3917 1384 3923 1396
rect 3933 1364 3939 1396
rect 4013 1344 4019 1476
rect 4045 1424 4051 1436
rect 4093 1364 4099 1436
rect 4109 1384 4115 1396
rect 3965 1244 3971 1316
rect 3981 1304 3987 1316
rect 4029 1244 4035 1316
rect 4077 1303 4083 1316
rect 4077 1297 4099 1303
rect 4093 1204 4099 1297
rect 3917 1184 3923 1196
rect 4125 1163 4131 1496
rect 4157 1424 4163 1496
rect 4173 1404 4179 1476
rect 4189 1464 4195 1497
rect 4205 1443 4211 1576
rect 4196 1437 4211 1443
rect 4141 1184 4147 1396
rect 4221 1384 4227 1676
rect 4173 1324 4179 1356
rect 4109 1157 4131 1163
rect 3892 1057 3900 1063
rect 3885 984 3891 1056
rect 3917 1004 3923 1116
rect 4045 1104 4051 1136
rect 3997 1044 4003 1096
rect 3917 984 3923 996
rect 3869 957 3891 963
rect 3741 926 3747 936
rect 3741 917 3747 918
rect 3828 917 3843 923
rect 3741 684 3747 796
rect 3821 784 3827 896
rect 3821 704 3827 756
rect 3709 483 3715 496
rect 3677 477 3715 483
rect 3709 424 3715 436
rect 3725 343 3731 676
rect 3741 604 3747 656
rect 3741 564 3747 596
rect 3757 584 3763 636
rect 3757 544 3763 556
rect 3773 544 3779 596
rect 3789 564 3795 596
rect 3805 544 3811 676
rect 3837 644 3843 917
rect 3860 897 3875 903
rect 3853 824 3859 856
rect 3853 704 3859 816
rect 3869 784 3875 897
rect 3885 804 3891 957
rect 3901 944 3907 956
rect 3981 944 3987 976
rect 4045 964 4051 1096
rect 4109 964 4115 1157
rect 4125 1064 4131 1136
rect 4173 1084 4179 1116
rect 3917 724 3923 816
rect 3917 704 3923 716
rect 3876 657 3891 663
rect 3837 564 3843 576
rect 3741 524 3747 536
rect 3780 517 3788 523
rect 3821 504 3827 556
rect 3853 544 3859 656
rect 3885 604 3891 657
rect 3869 504 3875 576
rect 3789 417 3843 423
rect 3789 364 3795 417
rect 3725 337 3747 343
rect 3524 297 3539 303
rect 3725 303 3731 316
rect 3668 297 3683 303
rect 3597 264 3603 276
rect 3565 184 3571 256
rect 3661 184 3667 236
rect 3677 203 3683 297
rect 3693 297 3731 303
rect 3693 284 3699 297
rect 3677 197 3699 203
rect 3693 184 3699 197
rect 3709 164 3715 196
rect 3524 117 3532 123
rect 3549 104 3555 156
rect 3725 144 3731 276
rect 3741 224 3747 337
rect 3764 297 3779 303
rect 3757 204 3763 276
rect 3773 243 3779 297
rect 3789 264 3795 336
rect 3805 304 3811 356
rect 3821 324 3827 396
rect 3837 324 3843 417
rect 3885 364 3891 596
rect 3901 424 3907 696
rect 3981 684 3987 936
rect 4157 924 4163 976
rect 3997 784 4003 816
rect 4029 724 4035 816
rect 4045 784 4051 918
rect 4141 844 4147 896
rect 4157 884 4163 916
rect 4173 763 4179 1076
rect 4205 1044 4211 1056
rect 4189 904 4195 956
rect 4221 924 4227 1096
rect 4237 943 4243 1696
rect 4253 1664 4259 1696
rect 4260 1617 4275 1623
rect 4269 1544 4275 1617
rect 4285 1504 4291 1716
rect 4301 1664 4307 1836
rect 4317 1804 4323 2076
rect 4349 2063 4355 2276
rect 4365 2124 4371 2256
rect 4381 2184 4387 2276
rect 4397 2104 4403 2396
rect 4429 2384 4435 2396
rect 4413 2324 4419 2336
rect 4445 2323 4451 2336
rect 4429 2317 4451 2323
rect 4429 2264 4435 2317
rect 4445 2244 4451 2296
rect 4461 2284 4467 2497
rect 4493 2483 4499 2577
rect 4509 2504 4515 2556
rect 4525 2524 4531 2716
rect 4589 2702 4595 2703
rect 4589 2684 4595 2694
rect 4541 2504 4547 2516
rect 4493 2477 4515 2483
rect 4477 2404 4483 2476
rect 4509 2384 4515 2477
rect 4525 2424 4531 2496
rect 4573 2444 4579 2536
rect 4621 2503 4627 2737
rect 4637 2524 4643 2836
rect 4664 2806 4665 2814
rect 4673 2806 4675 2814
rect 4683 2806 4685 2814
rect 4693 2806 4695 2814
rect 4703 2806 4712 2814
rect 4653 2664 4659 2696
rect 4765 2664 4771 2836
rect 4797 2704 4803 2716
rect 4845 2684 4851 2696
rect 4717 2584 4723 2636
rect 4765 2584 4771 2596
rect 4653 2564 4659 2576
rect 4861 2544 4867 2676
rect 4893 2664 4899 2676
rect 4877 2544 4883 2656
rect 4909 2644 4915 2676
rect 4973 2664 4979 2696
rect 4989 2540 4995 2576
rect 4733 2524 4739 2536
rect 4621 2497 4643 2503
rect 4477 2244 4483 2336
rect 4429 2124 4435 2176
rect 4477 2144 4483 2196
rect 4493 2164 4499 2316
rect 4509 2284 4515 2296
rect 4557 2204 4563 2236
rect 4445 2124 4451 2136
rect 4461 2124 4467 2136
rect 4413 2064 4419 2116
rect 4333 2057 4355 2063
rect 4333 1924 4339 2057
rect 4333 1763 4339 1876
rect 4381 1864 4387 1896
rect 4429 1864 4435 1976
rect 4445 1884 4451 2116
rect 4480 2096 4483 2103
rect 4365 1777 4419 1783
rect 4365 1764 4371 1777
rect 4413 1764 4419 1777
rect 4333 1757 4355 1763
rect 4324 1737 4332 1743
rect 4253 1404 4259 1496
rect 4269 1324 4275 1476
rect 4317 1384 4323 1556
rect 4349 1484 4355 1757
rect 4381 1664 4387 1756
rect 4365 1544 4371 1576
rect 4381 1544 4387 1656
rect 4397 1464 4403 1516
rect 4397 1444 4403 1456
rect 4413 1444 4419 1636
rect 4429 1544 4435 1736
rect 4477 1704 4483 2096
rect 4509 1964 4515 2056
rect 4573 1924 4579 2236
rect 4589 2164 4595 2196
rect 4589 2124 4595 2136
rect 4605 2064 4611 2196
rect 4621 2184 4627 2436
rect 4637 2284 4643 2497
rect 4749 2444 4755 2516
rect 4893 2504 4899 2518
rect 4925 2443 4931 2536
rect 5005 2503 5011 2536
rect 4989 2497 5011 2503
rect 4909 2437 4931 2443
rect 4664 2406 4665 2414
rect 4673 2406 4675 2414
rect 4683 2406 4685 2414
rect 4693 2406 4695 2414
rect 4703 2406 4712 2414
rect 4669 2304 4675 2376
rect 4653 2244 4659 2276
rect 4637 2184 4643 2236
rect 4749 2163 4755 2316
rect 4733 2157 4755 2163
rect 4701 2124 4707 2156
rect 4733 2144 4739 2157
rect 4605 1924 4611 1936
rect 4557 1844 4563 1876
rect 4573 1824 4579 1836
rect 4589 1804 4595 1856
rect 4525 1724 4531 1796
rect 4461 1464 4467 1596
rect 4301 1244 4307 1336
rect 4397 1324 4403 1356
rect 4253 1184 4259 1236
rect 4317 1144 4323 1276
rect 4333 1184 4339 1296
rect 4349 1244 4355 1316
rect 4413 1283 4419 1336
rect 4477 1304 4483 1318
rect 4413 1277 4435 1283
rect 4333 1103 4339 1116
rect 4381 1104 4387 1216
rect 4413 1164 4419 1236
rect 4333 1097 4348 1103
rect 4301 1064 4307 1096
rect 4429 1084 4435 1277
rect 4493 1244 4499 1596
rect 4573 1584 4579 1616
rect 4589 1563 4595 1616
rect 4557 1557 4595 1563
rect 4509 1344 4515 1496
rect 4525 1324 4531 1456
rect 4557 1404 4563 1557
rect 4237 937 4252 943
rect 4157 757 4179 763
rect 4109 744 4115 756
rect 4061 724 4067 736
rect 4029 704 4035 716
rect 4132 697 4147 703
rect 3917 623 3923 636
rect 3917 617 3939 623
rect 3917 524 3923 556
rect 3933 523 3939 617
rect 3981 584 3987 656
rect 4013 624 4019 696
rect 3997 604 4003 616
rect 3997 544 4003 596
rect 4013 524 4019 556
rect 4029 544 4035 636
rect 3933 517 3955 523
rect 3933 484 3939 496
rect 3869 304 3875 316
rect 3885 284 3891 356
rect 3901 324 3907 396
rect 3917 384 3923 436
rect 3933 384 3939 436
rect 3933 344 3939 376
rect 3917 284 3923 296
rect 3773 237 3795 243
rect 3773 144 3779 196
rect 3789 184 3795 237
rect 3805 164 3811 256
rect 3821 144 3827 156
rect 3645 104 3651 116
rect 3677 64 3683 116
rect 3773 104 3779 136
rect 3853 104 3859 136
rect 3885 124 3891 276
rect 3949 263 3955 517
rect 4093 523 4099 636
rect 4061 517 4099 523
rect 4061 504 4067 517
rect 3965 304 3971 456
rect 4061 384 4067 436
rect 4029 323 4035 356
rect 4029 317 4051 323
rect 3933 257 3955 263
rect 3901 124 3907 256
rect 3933 203 3939 257
rect 3965 224 3971 276
rect 3933 197 3955 203
rect 3949 183 3955 197
rect 3981 184 3987 216
rect 3949 177 3971 183
rect 3965 164 3971 177
rect 3917 144 3923 156
rect 3997 143 4003 236
rect 4029 224 4035 296
rect 4045 284 4051 317
rect 4109 304 4115 656
rect 4141 604 4147 697
rect 4157 684 4163 757
rect 4189 723 4195 876
rect 4205 744 4211 836
rect 4221 784 4227 896
rect 4237 884 4243 916
rect 4205 724 4211 736
rect 4173 717 4195 723
rect 4173 683 4179 717
rect 4205 684 4211 696
rect 4173 677 4188 683
rect 4157 644 4163 656
rect 4141 564 4147 596
rect 4157 584 4163 636
rect 4205 564 4211 676
rect 4221 663 4227 696
rect 4237 684 4243 716
rect 4253 684 4259 936
rect 4269 924 4275 976
rect 4317 924 4323 976
rect 4333 903 4339 1056
rect 4397 1043 4403 1056
rect 4397 1037 4435 1043
rect 4365 984 4371 1036
rect 4429 1023 4435 1037
rect 4461 1023 4467 1216
rect 4477 1044 4483 1096
rect 4429 1017 4483 1023
rect 4477 984 4483 1017
rect 4493 1003 4499 1236
rect 4509 1184 4515 1236
rect 4525 1184 4531 1316
rect 4541 1183 4547 1296
rect 4541 1177 4563 1183
rect 4525 1144 4531 1176
rect 4525 1104 4531 1136
rect 4557 1124 4563 1177
rect 4573 1063 4579 1376
rect 4605 1124 4611 1896
rect 4621 1423 4627 2116
rect 4637 2024 4643 2056
rect 4664 2006 4665 2014
rect 4673 2006 4675 2014
rect 4683 2006 4685 2014
rect 4693 2006 4695 2014
rect 4703 2006 4712 2014
rect 4733 1984 4739 2116
rect 4749 2084 4755 2116
rect 4765 2044 4771 2376
rect 4797 2244 4803 2256
rect 4861 2244 4867 2256
rect 4781 2184 4787 2196
rect 4797 2044 4803 2156
rect 4813 2024 4819 2176
rect 4861 2163 4867 2236
rect 4861 2157 4883 2163
rect 4877 2144 4883 2157
rect 4861 2124 4867 2136
rect 4877 2064 4883 2116
rect 4653 1804 4659 1896
rect 4685 1744 4691 1896
rect 4701 1784 4707 1976
rect 4845 1944 4851 2036
rect 4877 1963 4883 2056
rect 4909 1984 4915 2437
rect 4989 2324 4995 2497
rect 4925 2184 4931 2296
rect 4989 2144 4995 2316
rect 5037 2244 5043 2936
rect 5101 2723 5107 3236
rect 5405 3204 5411 3316
rect 5437 3284 5443 3316
rect 5472 3296 5475 3303
rect 5469 3284 5475 3296
rect 5517 3283 5523 3376
rect 5597 3364 5603 3476
rect 5645 3463 5651 3476
rect 5693 3463 5699 3477
rect 5645 3457 5699 3463
rect 5741 3444 5747 3476
rect 5773 3404 5779 3516
rect 5789 3503 5795 3596
rect 5805 3563 5811 3796
rect 5821 3744 5827 3776
rect 5821 3684 5827 3716
rect 5837 3644 5843 3736
rect 5853 3624 5859 3716
rect 5805 3557 5827 3563
rect 5805 3524 5811 3536
rect 5789 3497 5811 3503
rect 5549 3344 5555 3356
rect 5645 3343 5651 3356
rect 5629 3337 5651 3343
rect 5549 3303 5555 3336
rect 5613 3324 5619 3336
rect 5581 3304 5587 3316
rect 5549 3297 5564 3303
rect 5629 3303 5635 3337
rect 5661 3304 5667 3356
rect 5709 3324 5715 3356
rect 5741 3304 5747 3336
rect 5597 3297 5635 3303
rect 5597 3283 5603 3297
rect 5517 3277 5603 3283
rect 5757 3164 5763 3336
rect 5805 3304 5811 3497
rect 5821 3384 5827 3557
rect 5853 3523 5859 3576
rect 5869 3544 5875 3817
rect 5885 3784 5891 3877
rect 5933 3764 5939 3876
rect 5901 3724 5907 3736
rect 5885 3584 5891 3696
rect 5901 3563 5907 3656
rect 5917 3644 5923 3736
rect 5949 3723 5955 3916
rect 5965 3903 5971 3996
rect 5981 3924 5987 4036
rect 5997 3984 6003 4096
rect 6061 4084 6067 4116
rect 6093 4084 6099 4157
rect 6125 4144 6131 4176
rect 6141 4124 6147 4317
rect 6173 4304 6179 4356
rect 6221 4304 6227 4316
rect 6189 4224 6195 4256
rect 6125 4084 6131 4116
rect 5965 3897 5987 3903
rect 5965 3744 5971 3856
rect 5949 3717 5971 3723
rect 5885 3557 5907 3563
rect 5853 3517 5868 3523
rect 5837 3504 5843 3516
rect 5885 3504 5891 3557
rect 5933 3503 5939 3616
rect 5949 3584 5955 3696
rect 5965 3624 5971 3717
rect 5981 3624 5987 3897
rect 6013 3824 6019 3956
rect 6029 3904 6035 3976
rect 6061 3904 6067 4056
rect 6141 4024 6147 4096
rect 6157 4004 6163 4176
rect 6189 4144 6195 4156
rect 6221 4124 6227 4216
rect 6269 4144 6275 4256
rect 6173 4104 6179 4116
rect 6189 4104 6195 4116
rect 6173 3917 6211 3923
rect 6125 3904 6131 3916
rect 6173 3903 6179 3917
rect 6164 3897 6179 3903
rect 6109 3883 6115 3896
rect 6125 3884 6131 3896
rect 6205 3884 6211 3917
rect 6084 3877 6115 3883
rect 6148 3877 6163 3883
rect 5997 3784 6003 3796
rect 6029 3744 6035 3876
rect 6045 3824 6051 3876
rect 6061 3744 6067 3876
rect 6157 3864 6163 3877
rect 6157 3804 6163 3836
rect 6173 3824 6179 3876
rect 6189 3764 6195 3876
rect 6189 3744 6195 3756
rect 5917 3497 5939 3503
rect 5885 3484 5891 3496
rect 5917 3424 5923 3497
rect 5933 3464 5939 3476
rect 5949 3404 5955 3536
rect 5997 3524 6003 3696
rect 6013 3644 6019 3736
rect 6045 3704 6051 3716
rect 6093 3623 6099 3696
rect 6109 3684 6115 3736
rect 6125 3704 6131 3716
rect 6157 3704 6163 3716
rect 6205 3704 6211 3856
rect 6221 3804 6227 3916
rect 6237 3904 6243 4076
rect 6285 3944 6291 4096
rect 6253 3784 6259 3916
rect 6285 3844 6291 3936
rect 6077 3617 6099 3623
rect 6157 3623 6163 3696
rect 6157 3617 6179 3623
rect 5965 3464 5971 3476
rect 5821 3357 5859 3363
rect 5821 3344 5827 3357
rect 5837 3184 5843 3336
rect 5853 3324 5859 3357
rect 5876 3357 5907 3363
rect 5901 3344 5907 3357
rect 5901 3304 5907 3316
rect 5949 3284 5955 3316
rect 5981 3304 5987 3436
rect 5997 3364 6003 3396
rect 6013 3344 6019 3376
rect 6029 3344 6035 3616
rect 6077 3564 6083 3617
rect 6045 3464 6051 3516
rect 6077 3504 6083 3556
rect 6077 3444 6083 3456
rect 5165 2944 5171 3156
rect 5181 2984 5187 3116
rect 5197 3064 5203 3076
rect 5213 2944 5219 2956
rect 5149 2924 5155 2936
rect 5213 2904 5219 2916
rect 5117 2884 5123 2896
rect 5101 2717 5123 2723
rect 5117 2704 5123 2717
rect 5069 2664 5075 2676
rect 5069 2603 5075 2656
rect 5069 2597 5091 2603
rect 5085 2524 5091 2597
rect 5069 2364 5075 2396
rect 5005 2164 5011 2236
rect 5021 2184 5027 2196
rect 4877 1957 4899 1963
rect 4733 1884 4739 1936
rect 4829 1904 4835 1916
rect 4788 1897 4812 1903
rect 4749 1883 4755 1896
rect 4877 1884 4883 1936
rect 4893 1904 4899 1957
rect 4925 1924 4931 2116
rect 4749 1877 4764 1883
rect 4765 1844 4771 1856
rect 4701 1744 4707 1776
rect 4717 1724 4723 1796
rect 4765 1764 4771 1836
rect 4813 1824 4819 1856
rect 4861 1744 4867 1856
rect 4893 1784 4899 1816
rect 4909 1744 4915 1896
rect 4957 1823 4963 1916
rect 4989 1863 4995 1896
rect 5005 1884 5011 2136
rect 5037 2104 5043 2116
rect 5021 1884 5027 2016
rect 5037 1984 5043 2056
rect 5053 1944 5059 2136
rect 5069 2124 5075 2356
rect 5085 2284 5091 2516
rect 5101 2504 5107 2696
rect 5101 2304 5107 2496
rect 5117 2323 5123 2696
rect 5229 2684 5235 2996
rect 5261 2984 5267 2996
rect 5277 2924 5283 2936
rect 5293 2924 5299 3016
rect 5309 2944 5315 3116
rect 5325 3104 5331 3156
rect 5460 3117 5475 3123
rect 5469 3104 5475 3117
rect 5533 3084 5539 3116
rect 5373 2964 5379 3056
rect 5421 3043 5427 3076
rect 5453 3063 5459 3076
rect 5485 3063 5491 3076
rect 5453 3057 5491 3063
rect 5405 3037 5427 3043
rect 5389 2944 5395 3016
rect 5405 2984 5411 3037
rect 5437 2964 5443 3056
rect 5517 2964 5523 3076
rect 5533 3044 5539 3076
rect 5597 3064 5603 3116
rect 5629 3104 5635 3136
rect 5757 3084 5763 3156
rect 5796 3097 5827 3103
rect 5821 3083 5827 3097
rect 5821 3077 5843 3083
rect 5549 3057 5564 3063
rect 5549 3023 5555 3057
rect 5533 3017 5555 3023
rect 5421 2944 5427 2956
rect 5261 2724 5267 2896
rect 5325 2864 5331 2896
rect 5501 2864 5507 2956
rect 5517 2944 5523 2956
rect 5533 2924 5539 3017
rect 5517 2884 5523 2916
rect 5277 2784 5283 2856
rect 5277 2724 5283 2776
rect 5501 2744 5507 2836
rect 5264 2717 5267 2724
rect 5341 2702 5347 2716
rect 5309 2664 5315 2676
rect 5220 2657 5267 2663
rect 5261 2643 5267 2657
rect 5261 2637 5299 2643
rect 5293 2624 5299 2637
rect 5501 2624 5507 2636
rect 5341 2564 5347 2616
rect 5325 2544 5331 2556
rect 5389 2544 5395 2596
rect 5421 2557 5475 2563
rect 5133 2524 5139 2536
rect 5213 2504 5219 2516
rect 5229 2404 5235 2516
rect 5261 2384 5267 2416
rect 5117 2317 5139 2323
rect 5117 2283 5123 2296
rect 5101 2277 5123 2283
rect 5085 2144 5091 2156
rect 5101 2064 5107 2277
rect 5085 1924 5091 1936
rect 5069 1904 5075 1916
rect 5037 1863 5043 1896
rect 5085 1884 5091 1916
rect 5133 1904 5139 2317
rect 5213 2284 5219 2336
rect 5277 2304 5283 2536
rect 5421 2524 5427 2557
rect 5469 2543 5475 2557
rect 5469 2537 5484 2543
rect 5517 2543 5523 2736
rect 5549 2684 5555 2956
rect 5613 2924 5619 3036
rect 5629 2924 5635 2936
rect 5645 2924 5651 2956
rect 5661 2944 5667 3036
rect 5677 2984 5683 2996
rect 5693 2984 5699 3056
rect 5725 3044 5731 3056
rect 5741 2964 5747 3036
rect 5773 2984 5779 3076
rect 5789 3024 5795 3056
rect 5837 3044 5843 3077
rect 5581 2864 5587 2896
rect 5629 2804 5635 2916
rect 5677 2824 5683 2956
rect 5693 2904 5699 2936
rect 5709 2844 5715 2916
rect 5725 2864 5731 2936
rect 5741 2924 5747 2936
rect 5805 2924 5811 2976
rect 5757 2897 5772 2903
rect 5565 2704 5571 2716
rect 5597 2703 5603 2796
rect 5597 2697 5635 2703
rect 5629 2683 5635 2697
rect 5629 2677 5676 2683
rect 5709 2663 5715 2836
rect 5725 2764 5731 2856
rect 5757 2784 5763 2897
rect 5805 2764 5811 2836
rect 5725 2724 5731 2756
rect 5700 2657 5715 2663
rect 5549 2644 5555 2656
rect 5709 2604 5715 2636
rect 5741 2624 5747 2756
rect 5773 2723 5779 2736
rect 5773 2717 5811 2723
rect 5805 2704 5811 2717
rect 5789 2624 5795 2696
rect 5805 2664 5811 2676
rect 5501 2537 5523 2543
rect 5437 2524 5443 2536
rect 5501 2524 5507 2537
rect 5693 2524 5699 2536
rect 5437 2484 5443 2516
rect 5517 2504 5523 2516
rect 5629 2504 5635 2516
rect 5725 2504 5731 2536
rect 5757 2524 5763 2536
rect 5613 2444 5619 2496
rect 5725 2444 5731 2496
rect 5805 2484 5811 2516
rect 5597 2383 5603 2436
rect 5597 2377 5619 2383
rect 5613 2324 5619 2377
rect 5517 2284 5523 2296
rect 5677 2284 5683 2296
rect 5693 2284 5699 2436
rect 5165 2184 5171 2216
rect 5181 2164 5187 2176
rect 5213 2144 5219 2276
rect 5149 2104 5155 2116
rect 5204 2037 5219 2043
rect 5213 1944 5219 2037
rect 5229 1944 5235 2236
rect 5261 2124 5267 2236
rect 5517 2164 5523 2276
rect 5677 2164 5683 2196
rect 5325 2064 5331 2076
rect 5325 1944 5331 2056
rect 5197 1924 5203 1936
rect 5341 1924 5347 1936
rect 5357 1924 5363 2116
rect 5405 1924 5411 1936
rect 5357 1917 5360 1924
rect 5421 1904 5427 2116
rect 5501 1944 5507 2136
rect 4989 1857 5011 1863
rect 5037 1857 5084 1863
rect 4941 1817 4963 1823
rect 4941 1784 4947 1817
rect 5005 1784 5011 1857
rect 5117 1824 5123 1896
rect 5133 1864 5139 1876
rect 5117 1784 5123 1816
rect 4989 1764 4995 1776
rect 4797 1704 4803 1716
rect 4813 1664 4819 1696
rect 4861 1644 4867 1716
rect 4884 1697 4899 1703
rect 4845 1624 4851 1636
rect 4664 1606 4665 1614
rect 4673 1606 4675 1614
rect 4683 1606 4685 1614
rect 4693 1606 4695 1614
rect 4703 1606 4712 1614
rect 4637 1544 4643 1596
rect 4669 1544 4675 1576
rect 4685 1524 4691 1576
rect 4733 1544 4739 1596
rect 4877 1584 4883 1656
rect 4733 1484 4739 1516
rect 4813 1484 4819 1496
rect 4829 1484 4835 1516
rect 4621 1417 4643 1423
rect 4621 1384 4627 1396
rect 4573 1057 4595 1063
rect 4589 1044 4595 1057
rect 4493 997 4515 1003
rect 4493 943 4499 976
rect 4477 937 4499 943
rect 4413 904 4419 936
rect 4477 904 4483 937
rect 4509 924 4515 997
rect 4541 923 4547 1016
rect 4605 944 4611 976
rect 4637 924 4643 1417
rect 4653 1344 4659 1396
rect 4669 1384 4675 1456
rect 4717 1284 4723 1436
rect 4781 1404 4787 1436
rect 4829 1344 4835 1396
rect 4845 1384 4851 1456
rect 4861 1444 4867 1536
rect 4877 1504 4883 1516
rect 4893 1483 4899 1697
rect 4925 1684 4931 1756
rect 5069 1744 5075 1756
rect 4909 1584 4915 1656
rect 4957 1624 4963 1736
rect 4973 1724 4979 1736
rect 5021 1703 5027 1736
rect 5037 1724 5043 1736
rect 5021 1697 5043 1703
rect 4941 1484 4947 1496
rect 4877 1477 4899 1483
rect 4664 1206 4665 1214
rect 4673 1206 4675 1214
rect 4683 1206 4685 1214
rect 4693 1206 4695 1214
rect 4703 1206 4712 1214
rect 4733 1184 4739 1336
rect 4653 1104 4659 1116
rect 4541 917 4563 923
rect 4333 897 4348 903
rect 4509 903 4515 916
rect 4500 897 4515 903
rect 4557 903 4563 917
rect 4557 897 4579 903
rect 4285 743 4291 876
rect 4285 737 4307 743
rect 4301 724 4307 737
rect 4269 684 4275 696
rect 4333 683 4339 796
rect 4349 743 4355 876
rect 4365 824 4371 896
rect 4349 737 4371 743
rect 4365 724 4371 737
rect 4349 704 4355 716
rect 4381 704 4387 796
rect 4365 697 4380 703
rect 4365 684 4371 697
rect 4333 677 4355 683
rect 4221 657 4243 663
rect 4237 584 4243 657
rect 4125 524 4131 536
rect 4205 524 4211 536
rect 4141 484 4147 516
rect 4068 297 4083 303
rect 4077 243 4083 297
rect 4109 284 4115 296
rect 4157 284 4163 356
rect 4173 304 4179 356
rect 4189 344 4195 516
rect 4253 504 4259 516
rect 4269 484 4275 616
rect 4301 584 4307 636
rect 4317 564 4323 636
rect 4285 484 4291 556
rect 4221 384 4227 396
rect 4141 244 4147 256
rect 4045 237 4083 243
rect 4045 203 4051 237
rect 3981 137 4003 143
rect 4013 197 4051 203
rect 3901 104 3907 116
rect 3876 97 3884 103
rect 3965 63 3971 116
rect 3981 84 3987 137
rect 4013 123 4019 197
rect 4141 164 4147 176
rect 4109 124 4115 136
rect 3997 117 4019 123
rect 3997 63 4003 117
rect 4061 117 4076 123
rect 4045 104 4051 116
rect 4061 104 4067 117
rect 4084 97 4092 103
rect 4125 84 4131 116
rect 4189 104 4195 156
rect 3965 57 4003 63
rect 4205 44 4211 376
rect 4221 163 4227 176
rect 4237 163 4243 376
rect 4285 164 4291 476
rect 4317 443 4323 516
rect 4333 504 4339 536
rect 4349 524 4355 677
rect 4317 437 4339 443
rect 4317 303 4323 416
rect 4333 364 4339 437
rect 4365 323 4371 436
rect 4397 424 4403 896
rect 4541 884 4547 896
rect 4413 703 4419 816
rect 4429 724 4435 876
rect 4573 863 4579 897
rect 4461 857 4499 863
rect 4573 857 4611 863
rect 4461 823 4467 857
rect 4445 817 4467 823
rect 4445 784 4451 817
rect 4493 804 4499 857
rect 4509 824 4515 836
rect 4573 824 4579 836
rect 4525 817 4563 823
rect 4461 763 4467 796
rect 4461 757 4483 763
rect 4477 724 4483 757
rect 4509 723 4515 816
rect 4525 804 4531 817
rect 4557 763 4563 817
rect 4589 784 4595 836
rect 4605 763 4611 857
rect 4621 784 4627 896
rect 4557 757 4595 763
rect 4605 757 4627 763
rect 4509 717 4563 723
rect 4413 697 4428 703
rect 4461 703 4467 716
rect 4493 704 4499 716
rect 4461 697 4483 703
rect 4477 683 4483 697
rect 4557 703 4563 717
rect 4589 703 4595 757
rect 4621 724 4627 757
rect 4637 723 4643 896
rect 4669 884 4675 1156
rect 4749 1143 4755 1336
rect 4765 1304 4771 1316
rect 4733 1137 4755 1143
rect 4733 1124 4739 1137
rect 4733 1104 4739 1116
rect 4781 1084 4787 1216
rect 4797 1124 4803 1136
rect 4829 1104 4835 1176
rect 4845 1104 4851 1316
rect 4861 1304 4867 1376
rect 4877 1144 4883 1477
rect 4909 1444 4915 1476
rect 4893 1324 4899 1416
rect 4909 1344 4915 1436
rect 4989 1404 4995 1476
rect 5005 1464 5011 1636
rect 5021 1504 5027 1536
rect 5037 1484 5043 1697
rect 5069 1644 5075 1716
rect 5069 1504 5075 1636
rect 5085 1624 5091 1736
rect 5117 1723 5123 1776
rect 5133 1744 5139 1856
rect 5245 1824 5251 1896
rect 5316 1877 5324 1883
rect 5261 1864 5267 1876
rect 5453 1864 5459 1876
rect 5245 1757 5283 1763
rect 5117 1717 5132 1723
rect 5149 1664 5155 1736
rect 5245 1704 5251 1757
rect 5277 1723 5283 1757
rect 5437 1744 5443 1776
rect 5469 1764 5475 1836
rect 5501 1824 5507 1856
rect 5485 1724 5491 1816
rect 5533 1784 5539 1876
rect 5277 1717 5299 1723
rect 5085 1584 5091 1616
rect 4957 1324 4963 1356
rect 4909 1317 4947 1323
rect 4909 1184 4915 1317
rect 4941 1304 4947 1317
rect 4973 1323 4979 1336
rect 4973 1317 4995 1323
rect 4973 1184 4979 1236
rect 4925 1157 4963 1163
rect 4685 963 4691 1076
rect 4701 1024 4707 1036
rect 4781 984 4787 1016
rect 4685 957 4755 963
rect 4749 944 4755 957
rect 4717 843 4723 936
rect 4717 837 4739 843
rect 4664 806 4665 814
rect 4673 806 4675 814
rect 4683 806 4685 814
rect 4693 806 4695 814
rect 4703 806 4712 814
rect 4637 717 4659 723
rect 4557 697 4579 703
rect 4589 697 4636 703
rect 4525 683 4531 696
rect 4477 677 4531 683
rect 4573 664 4579 697
rect 4413 623 4419 656
rect 4445 637 4460 643
rect 4413 617 4435 623
rect 4413 524 4419 596
rect 4429 463 4435 617
rect 4445 484 4451 637
rect 4461 524 4467 616
rect 4493 603 4499 656
rect 4477 597 4499 603
rect 4429 457 4451 463
rect 4429 344 4435 436
rect 4349 317 4371 323
rect 4317 297 4339 303
rect 4301 284 4307 296
rect 4333 284 4339 297
rect 4317 263 4323 276
rect 4349 263 4355 317
rect 4365 297 4412 303
rect 4365 284 4371 297
rect 4317 257 4355 263
rect 4221 157 4243 163
rect 4221 124 4227 157
rect 4237 104 4243 136
rect 4269 103 4275 156
rect 4285 144 4291 156
rect 4317 124 4323 257
rect 4333 184 4339 236
rect 4349 163 4355 236
rect 4381 224 4387 276
rect 4429 264 4435 316
rect 4333 157 4355 163
rect 4253 97 4275 103
rect 4221 83 4227 96
rect 4253 83 4259 97
rect 4221 77 4259 83
rect 4333 64 4339 157
rect 4445 163 4451 457
rect 4477 404 4483 597
rect 4493 524 4499 576
rect 4525 504 4531 636
rect 4589 583 4595 636
rect 4637 603 4643 676
rect 4653 644 4659 717
rect 4669 684 4675 776
rect 4733 744 4739 837
rect 4717 703 4723 736
rect 4749 704 4755 816
rect 4765 744 4771 876
rect 4765 724 4771 736
rect 4692 697 4723 703
rect 4797 683 4803 1036
rect 4813 963 4819 1096
rect 4845 1044 4851 1076
rect 4909 1023 4915 1136
rect 4925 1104 4931 1157
rect 4941 1124 4947 1136
rect 4941 1083 4947 1116
rect 4932 1077 4947 1083
rect 4957 1063 4963 1157
rect 4989 1104 4995 1317
rect 5037 1264 5043 1476
rect 5053 1424 5059 1436
rect 5021 1184 5027 1256
rect 5005 1103 5011 1136
rect 5053 1124 5059 1356
rect 5101 1324 5107 1416
rect 5149 1403 5155 1656
rect 5261 1564 5267 1716
rect 5293 1704 5299 1717
rect 5389 1704 5395 1716
rect 5517 1704 5523 1756
rect 5533 1704 5539 1756
rect 5549 1744 5555 1896
rect 5277 1684 5283 1696
rect 5277 1524 5283 1616
rect 5293 1537 5331 1543
rect 5293 1524 5299 1537
rect 5213 1502 5219 1516
rect 5325 1504 5331 1537
rect 5245 1484 5251 1496
rect 5245 1464 5251 1476
rect 5133 1397 5155 1403
rect 5133 1364 5139 1397
rect 5165 1377 5180 1383
rect 5165 1364 5171 1377
rect 5069 1224 5075 1256
rect 5085 1244 5091 1316
rect 5092 1237 5100 1243
rect 5005 1097 5027 1103
rect 5021 1083 5027 1097
rect 5021 1077 5043 1083
rect 4861 1017 4915 1023
rect 4941 1057 4963 1063
rect 4813 957 4851 963
rect 4829 784 4835 936
rect 4829 764 4835 776
rect 4829 704 4835 716
rect 4845 704 4851 957
rect 4861 784 4867 1017
rect 4893 997 4931 1003
rect 4893 984 4899 997
rect 4925 984 4931 997
rect 4893 924 4899 956
rect 4909 903 4915 976
rect 4941 963 4947 1057
rect 4973 1043 4979 1076
rect 4989 1044 4995 1076
rect 5005 1064 5011 1076
rect 5037 1063 5043 1077
rect 5069 1083 5075 1216
rect 5133 1164 5139 1296
rect 5149 1184 5155 1216
rect 5133 1144 5139 1156
rect 5101 1104 5107 1136
rect 5117 1084 5123 1116
rect 5149 1084 5155 1096
rect 5060 1077 5075 1083
rect 5181 1083 5187 1116
rect 5165 1077 5187 1083
rect 5037 1057 5139 1063
rect 4932 957 4947 963
rect 4957 1037 4979 1043
rect 4893 897 4915 903
rect 4893 884 4899 897
rect 4909 784 4915 876
rect 4941 823 4947 896
rect 4957 884 4963 1037
rect 4973 943 4979 1016
rect 4989 997 5027 1003
rect 4989 984 4995 997
rect 5021 984 5027 997
rect 4973 937 4988 943
rect 4925 817 4947 823
rect 4925 704 4931 817
rect 4941 724 4947 756
rect 4797 677 4835 683
rect 4557 577 4595 583
rect 4621 597 4643 603
rect 4493 484 4499 496
rect 4493 404 4499 476
rect 4525 384 4531 396
rect 4541 363 4547 516
rect 4557 404 4563 577
rect 4621 563 4627 597
rect 4596 557 4627 563
rect 4653 544 4659 576
rect 4621 523 4627 536
rect 4605 517 4627 523
rect 4477 357 4547 363
rect 4461 284 4467 356
rect 4477 324 4483 357
rect 4493 304 4499 336
rect 4509 324 4515 336
rect 4541 324 4547 336
rect 4557 304 4563 356
rect 4477 283 4483 296
rect 4589 284 4595 456
rect 4605 404 4611 517
rect 4685 444 4691 636
rect 4717 623 4723 656
rect 4765 644 4771 676
rect 4813 643 4819 656
rect 4797 637 4819 643
rect 4701 617 4723 623
rect 4701 523 4707 617
rect 4701 517 4723 523
rect 4701 464 4707 496
rect 4717 443 4723 517
rect 4717 437 4739 443
rect 4605 344 4611 376
rect 4477 277 4515 283
rect 4509 263 4515 277
rect 4509 257 4556 263
rect 4461 244 4467 256
rect 4493 243 4499 256
rect 4605 244 4611 296
rect 4621 284 4627 356
rect 4637 323 4643 436
rect 4664 406 4665 414
rect 4673 406 4675 414
rect 4683 406 4685 414
rect 4693 406 4695 414
rect 4703 406 4712 414
rect 4733 404 4739 437
rect 4733 344 4739 396
rect 4637 317 4684 323
rect 4749 323 4755 376
rect 4765 363 4771 636
rect 4797 584 4803 637
rect 4797 543 4803 576
rect 4781 537 4803 543
rect 4781 524 4787 537
rect 4797 503 4803 516
rect 4829 504 4835 677
rect 4877 624 4883 656
rect 4925 644 4931 656
rect 4957 644 4963 796
rect 4973 724 4979 916
rect 5005 704 5011 756
rect 5021 724 5027 876
rect 5037 704 5043 1016
rect 5053 924 5059 1036
rect 5069 884 5075 896
rect 5069 824 5075 836
rect 5085 824 5091 1016
rect 5133 984 5139 1057
rect 5101 924 5107 936
rect 5117 884 5123 956
rect 5149 924 5155 956
rect 5069 784 5075 816
rect 5101 784 5107 876
rect 5133 764 5139 816
rect 5149 784 5155 816
rect 5165 764 5171 1077
rect 5181 924 5187 1036
rect 5197 944 5203 1356
rect 5293 1344 5299 1456
rect 5309 1424 5315 1496
rect 5325 1464 5331 1476
rect 5405 1464 5411 1476
rect 5277 1324 5283 1336
rect 5309 1284 5315 1316
rect 5213 1224 5219 1276
rect 5213 1104 5219 1216
rect 5293 1144 5299 1276
rect 5341 1244 5347 1356
rect 5421 1344 5427 1456
rect 5309 1184 5315 1216
rect 5293 1123 5299 1136
rect 5341 1124 5347 1156
rect 5293 1117 5315 1123
rect 5277 1103 5283 1116
rect 5277 1097 5292 1103
rect 5309 1103 5315 1117
rect 5373 1104 5379 1116
rect 5309 1097 5331 1103
rect 5325 1084 5331 1097
rect 5245 1044 5251 1056
rect 5309 1044 5315 1076
rect 5389 1063 5395 1076
rect 5373 1057 5395 1063
rect 5325 1044 5331 1056
rect 5373 1044 5379 1057
rect 5405 1044 5411 1256
rect 5437 1104 5443 1676
rect 5453 1584 5459 1656
rect 5565 1644 5571 1936
rect 5581 1924 5587 2036
rect 5597 1944 5603 2136
rect 5677 2124 5683 2136
rect 5613 2024 5619 2036
rect 5613 1784 5619 1816
rect 5661 1784 5667 1916
rect 5693 1863 5699 2256
rect 5709 2204 5715 2276
rect 5709 1904 5715 1976
rect 5725 1864 5731 2416
rect 5741 2324 5747 2436
rect 5741 2304 5747 2316
rect 5757 2203 5763 2236
rect 5741 2197 5763 2203
rect 5741 2126 5747 2197
rect 5741 2117 5747 2118
rect 5773 2024 5779 2376
rect 5821 2304 5827 2636
rect 5837 2544 5843 3036
rect 5869 3004 5875 3256
rect 5901 3164 5907 3236
rect 5949 3184 5955 3236
rect 5949 3124 5955 3176
rect 5901 3103 5907 3116
rect 5885 3097 5907 3103
rect 5885 3084 5891 3097
rect 5917 3037 5948 3043
rect 5917 3003 5923 3037
rect 5901 2997 5923 3003
rect 5869 2824 5875 2996
rect 5885 2864 5891 2916
rect 5901 2904 5907 2997
rect 5965 2964 5971 3156
rect 5981 3144 5987 3296
rect 5997 3164 6003 3236
rect 5981 3104 5987 3116
rect 6013 3103 6019 3316
rect 6029 3264 6035 3316
rect 6045 3264 6051 3416
rect 6061 3404 6067 3436
rect 6093 3424 6099 3596
rect 6173 3584 6179 3617
rect 6189 3504 6195 3696
rect 6205 3483 6211 3516
rect 6189 3477 6211 3483
rect 6189 3464 6195 3477
rect 6125 3444 6131 3456
rect 6141 3344 6147 3356
rect 6109 3303 6115 3316
rect 6141 3304 6147 3316
rect 6109 3297 6131 3303
rect 5997 3097 6019 3103
rect 5981 3064 5987 3076
rect 5965 2923 5971 2956
rect 5981 2944 5987 2956
rect 5965 2917 5980 2923
rect 5997 2904 6003 3097
rect 6029 3084 6035 3156
rect 5853 2704 5859 2776
rect 5885 2764 5891 2836
rect 5901 2724 5907 2736
rect 5904 2717 5907 2724
rect 5869 2704 5875 2716
rect 5917 2683 5923 2716
rect 5933 2704 5939 2716
rect 5917 2677 5932 2683
rect 5853 2624 5859 2676
rect 5933 2644 5939 2676
rect 5901 2424 5907 2616
rect 5949 2603 5955 2716
rect 5965 2644 5971 2896
rect 6013 2884 6019 3036
rect 6029 3003 6035 3076
rect 6045 3064 6051 3176
rect 6061 3124 6067 3296
rect 6125 3283 6131 3297
rect 6125 3277 6147 3283
rect 6093 3184 6099 3236
rect 6109 3083 6115 3256
rect 6093 3077 6115 3083
rect 6077 3064 6083 3076
rect 6029 2997 6051 3003
rect 6045 2944 6051 2997
rect 6029 2864 6035 2896
rect 5981 2724 5987 2736
rect 5997 2624 6003 2856
rect 6013 2784 6019 2796
rect 6013 2697 6051 2703
rect 6013 2664 6019 2697
rect 6029 2664 6035 2676
rect 6045 2664 6051 2697
rect 5949 2597 5971 2603
rect 5965 2544 5971 2597
rect 6013 2584 6019 2596
rect 5917 2504 5923 2516
rect 5933 2464 5939 2536
rect 5805 2284 5811 2296
rect 5940 2277 5948 2283
rect 5805 2124 5811 2236
rect 5821 2204 5827 2276
rect 5853 2164 5859 2236
rect 5821 2124 5827 2156
rect 5869 2124 5875 2196
rect 5949 2183 5955 2236
rect 5933 2177 5955 2183
rect 5933 2156 5939 2177
rect 5805 1984 5811 2116
rect 5917 2084 5923 2096
rect 5741 1864 5747 1956
rect 5821 1904 5827 1916
rect 5677 1857 5699 1863
rect 5581 1744 5587 1756
rect 5581 1664 5587 1716
rect 5597 1704 5603 1756
rect 5645 1744 5651 1776
rect 5629 1724 5635 1736
rect 5597 1684 5603 1696
rect 5613 1664 5619 1696
rect 5453 1324 5459 1416
rect 5485 1304 5491 1476
rect 5501 1384 5507 1516
rect 5549 1504 5555 1516
rect 5533 1344 5539 1496
rect 5549 1344 5555 1476
rect 5597 1383 5603 1636
rect 5629 1384 5635 1716
rect 5661 1704 5667 1716
rect 5677 1703 5683 1857
rect 5725 1783 5731 1836
rect 5709 1777 5731 1783
rect 5709 1744 5715 1777
rect 5789 1744 5795 1776
rect 5869 1764 5875 1796
rect 5677 1697 5699 1703
rect 5661 1504 5667 1576
rect 5597 1377 5612 1383
rect 5517 1184 5523 1196
rect 5277 1004 5283 1036
rect 5309 1023 5315 1036
rect 5309 1017 5347 1023
rect 5341 1003 5347 1017
rect 5341 997 5363 1003
rect 5357 984 5363 997
rect 5325 957 5356 963
rect 5325 944 5331 957
rect 5213 937 5228 943
rect 5213 924 5219 937
rect 5197 897 5212 903
rect 4973 643 4979 656
rect 4973 637 5011 643
rect 4941 583 4947 616
rect 4941 577 4963 583
rect 4877 544 4883 556
rect 4909 523 4915 576
rect 4925 544 4931 576
rect 4909 517 4924 523
rect 4788 497 4803 503
rect 4893 497 4924 503
rect 4781 383 4787 496
rect 4861 483 4867 496
rect 4861 477 4883 483
rect 4861 404 4867 436
rect 4804 397 4835 403
rect 4829 384 4835 397
rect 4781 377 4803 383
rect 4765 357 4787 363
rect 4733 317 4755 323
rect 4644 257 4659 263
rect 4493 237 4515 243
rect 4461 184 4467 236
rect 4445 157 4476 163
rect 4509 163 4515 237
rect 4509 157 4524 163
rect 4349 103 4355 136
rect 4365 124 4371 156
rect 4413 124 4419 156
rect 4461 137 4476 143
rect 4445 124 4451 136
rect 4381 104 4387 116
rect 4349 97 4371 103
rect 4365 83 4371 97
rect 4461 103 4467 137
rect 4493 104 4499 116
rect 4413 97 4467 103
rect 4365 77 4403 83
rect 4397 43 4403 77
rect 4413 64 4419 97
rect 4525 43 4531 116
rect 4541 64 4547 156
rect 4557 103 4563 176
rect 4589 163 4595 216
rect 4605 184 4611 196
rect 4621 164 4627 176
rect 4589 157 4611 163
rect 4605 103 4611 157
rect 4621 124 4627 156
rect 4637 103 4643 236
rect 4653 183 4659 257
rect 4669 204 4675 296
rect 4685 224 4691 276
rect 4653 177 4675 183
rect 4557 97 4595 103
rect 4605 97 4643 103
rect 4589 83 4595 97
rect 4589 77 4652 83
rect 4669 44 4675 177
rect 4397 37 4531 43
rect 4637 -17 4643 16
rect 4664 6 4665 14
rect 4673 6 4675 14
rect 4683 6 4685 14
rect 4693 6 4695 14
rect 4703 6 4712 14
rect 4733 -17 4739 317
rect 4749 244 4755 296
rect 4765 284 4771 336
rect 4781 263 4787 357
rect 4797 304 4803 377
rect 4813 304 4819 316
rect 4765 257 4787 263
rect 4765 224 4771 257
rect 4781 224 4787 236
rect 4797 164 4803 296
rect 4813 204 4819 276
rect 4829 144 4835 296
rect 4845 284 4851 356
rect 4877 304 4883 477
rect 4893 424 4899 497
rect 4909 463 4915 476
rect 4909 457 4931 463
rect 4925 324 4931 457
rect 4861 164 4867 276
rect 4877 224 4883 256
rect 4877 184 4883 196
rect 4861 124 4867 156
rect 4804 117 4812 123
rect 4781 103 4787 116
rect 4829 103 4835 116
rect 4781 97 4835 103
rect 4909 24 4915 296
rect 4925 124 4931 236
rect 4941 124 4947 456
rect 4957 404 4963 577
rect 4989 524 4995 596
rect 5005 584 5011 637
rect 5021 524 5027 636
rect 4957 264 4963 296
rect 4989 283 4995 496
rect 5037 484 5043 596
rect 5053 584 5059 636
rect 5069 543 5075 756
rect 5101 564 5107 756
rect 5156 717 5171 723
rect 5117 604 5123 676
rect 5149 664 5155 676
rect 5108 557 5123 563
rect 5117 543 5123 557
rect 5165 543 5171 717
rect 5197 584 5203 897
rect 5229 784 5235 916
rect 5245 664 5251 696
rect 5229 624 5235 636
rect 5213 544 5219 596
rect 5069 537 5107 543
rect 5117 537 5139 543
rect 5165 537 5187 543
rect 5076 517 5084 523
rect 5021 443 5027 456
rect 5021 437 5043 443
rect 5037 424 5043 437
rect 5069 364 5075 436
rect 5101 384 5107 537
rect 5133 464 5139 537
rect 5181 524 5187 537
rect 5149 363 5155 396
rect 5165 384 5171 516
rect 5133 357 5155 363
rect 5053 324 5059 336
rect 5021 284 5027 296
rect 4980 277 4995 283
rect 5085 263 5091 356
rect 5101 284 5107 296
rect 5117 264 5123 316
rect 5028 257 5075 263
rect 5085 257 5107 263
rect 5069 243 5075 257
rect 5069 237 5091 243
rect 4973 144 4979 216
rect 5037 164 5043 216
rect 5053 164 5059 236
rect 5085 184 5091 237
rect 5021 137 5068 143
rect 5021 123 5027 137
rect 5101 124 5107 257
rect 5133 184 5139 357
rect 5181 324 5187 516
rect 5213 484 5219 516
rect 5229 484 5235 556
rect 5245 543 5251 636
rect 5261 624 5267 896
rect 5277 784 5283 896
rect 5309 824 5315 916
rect 5341 903 5347 936
rect 5357 924 5363 956
rect 5341 897 5356 903
rect 5373 883 5379 1036
rect 5421 1004 5427 1076
rect 5437 964 5443 996
rect 5469 984 5475 1096
rect 5485 1064 5491 1136
rect 5549 1084 5555 1336
rect 5565 1164 5571 1296
rect 5581 1184 5587 1236
rect 5597 1204 5603 1336
rect 5485 1023 5491 1036
rect 5485 1017 5516 1023
rect 5389 943 5395 956
rect 5517 944 5523 996
rect 5533 984 5539 1076
rect 5565 1043 5571 1156
rect 5645 1143 5651 1436
rect 5677 1424 5683 1496
rect 5677 1324 5683 1336
rect 5693 1264 5699 1697
rect 5709 1344 5715 1676
rect 5725 1504 5731 1716
rect 5757 1564 5763 1716
rect 5869 1704 5875 1756
rect 5805 1664 5811 1696
rect 5837 1564 5843 1596
rect 5764 1517 5772 1523
rect 5725 1464 5731 1476
rect 5757 1403 5763 1476
rect 5741 1397 5763 1403
rect 5725 1304 5731 1316
rect 5725 1184 5731 1276
rect 5741 1163 5747 1397
rect 5741 1157 5763 1163
rect 5629 1137 5651 1143
rect 5597 1104 5603 1136
rect 5629 1104 5635 1137
rect 5549 1037 5571 1043
rect 5389 937 5404 943
rect 5341 877 5379 883
rect 5277 684 5283 756
rect 5325 704 5331 876
rect 5341 763 5347 877
rect 5364 777 5372 783
rect 5341 757 5363 763
rect 5357 723 5363 757
rect 5357 717 5388 723
rect 5300 677 5331 683
rect 5293 623 5299 656
rect 5277 617 5299 623
rect 5325 623 5331 677
rect 5357 644 5363 717
rect 5373 624 5379 696
rect 5421 664 5427 936
rect 5437 904 5443 936
rect 5533 924 5539 956
rect 5453 903 5459 916
rect 5453 897 5491 903
rect 5485 884 5491 897
rect 5437 864 5443 876
rect 5437 824 5443 856
rect 5453 803 5459 856
rect 5437 797 5459 803
rect 5469 803 5475 876
rect 5469 797 5491 803
rect 5325 617 5363 623
rect 5245 537 5267 543
rect 5149 184 5155 256
rect 5165 184 5171 256
rect 5197 244 5203 296
rect 5213 284 5219 316
rect 5229 264 5235 456
rect 5245 323 5251 516
rect 5261 364 5267 537
rect 5277 464 5283 617
rect 5341 484 5347 596
rect 5357 564 5363 617
rect 5421 584 5427 636
rect 5341 424 5347 436
rect 5245 317 5283 323
rect 5245 297 5260 303
rect 5213 257 5228 263
rect 5213 223 5219 257
rect 5245 244 5251 297
rect 5277 263 5283 317
rect 5277 257 5308 263
rect 5181 217 5219 223
rect 5181 184 5187 217
rect 5005 117 5027 123
rect 5005 103 5011 117
rect 5085 103 5091 116
rect 4948 97 5011 103
rect 5069 97 5091 103
rect 4941 84 4947 96
rect 5069 84 5075 97
rect 5117 63 5123 136
rect 5133 104 5139 136
rect 5213 64 5219 196
rect 5229 124 5235 236
rect 5261 84 5267 256
rect 5277 164 5283 236
rect 5325 184 5331 316
rect 5341 304 5347 416
rect 5357 304 5363 336
rect 5277 124 5283 156
rect 5341 144 5347 216
rect 5357 143 5363 296
rect 5373 164 5379 316
rect 5389 304 5395 496
rect 5421 484 5427 516
rect 5437 504 5443 797
rect 5469 764 5475 776
rect 5485 744 5491 797
rect 5501 704 5507 916
rect 5549 904 5555 1037
rect 5565 984 5571 1016
rect 5581 964 5587 1096
rect 5597 1023 5603 1076
rect 5613 1044 5619 1076
rect 5629 1023 5635 1036
rect 5597 1017 5635 1023
rect 5613 964 5619 996
rect 5597 924 5603 936
rect 5572 897 5603 903
rect 5517 684 5523 856
rect 5549 724 5555 876
rect 5565 684 5571 856
rect 5597 784 5603 897
rect 5613 864 5619 936
rect 5645 924 5651 1116
rect 5661 964 5667 1096
rect 5677 943 5683 1156
rect 5693 1117 5731 1123
rect 5693 1104 5699 1117
rect 5725 1104 5731 1117
rect 5709 964 5715 1076
rect 5725 1024 5731 1076
rect 5725 944 5731 1016
rect 5741 1003 5747 1136
rect 5757 1124 5763 1157
rect 5773 1144 5779 1476
rect 5789 1464 5795 1476
rect 5805 1384 5811 1396
rect 5773 1103 5779 1136
rect 5805 1104 5811 1316
rect 5821 1224 5827 1556
rect 5837 1524 5843 1556
rect 5837 1484 5843 1496
rect 5837 1183 5843 1376
rect 5869 1204 5875 1636
rect 5901 1623 5907 1836
rect 5885 1617 5907 1623
rect 5837 1177 5859 1183
rect 5837 1124 5843 1136
rect 5757 1097 5779 1103
rect 5757 1064 5763 1097
rect 5821 1084 5827 1116
rect 5741 997 5763 1003
rect 5757 984 5763 997
rect 5773 963 5779 1036
rect 5757 957 5779 963
rect 5677 937 5699 943
rect 5629 864 5635 896
rect 5597 703 5603 776
rect 5613 704 5619 776
rect 5629 704 5635 836
rect 5661 823 5667 856
rect 5677 844 5683 916
rect 5693 844 5699 937
rect 5757 943 5763 957
rect 5805 944 5811 1076
rect 5741 937 5763 943
rect 5661 817 5683 823
rect 5588 697 5603 703
rect 5645 684 5651 816
rect 5453 424 5459 656
rect 5469 624 5475 676
rect 5549 624 5555 676
rect 5565 604 5571 656
rect 5677 644 5683 817
rect 5709 784 5715 936
rect 5725 804 5731 916
rect 5741 884 5747 937
rect 5789 904 5795 916
rect 5805 764 5811 816
rect 5741 704 5747 756
rect 5773 717 5788 723
rect 5693 664 5699 696
rect 5492 557 5507 563
rect 5501 523 5507 557
rect 5485 517 5507 523
rect 5469 364 5475 496
rect 5485 404 5491 517
rect 5501 424 5507 476
rect 5517 404 5523 556
rect 5581 544 5587 636
rect 5597 523 5603 636
rect 5629 524 5635 616
rect 5645 584 5651 636
rect 5677 544 5683 596
rect 5709 544 5715 656
rect 5757 644 5763 656
rect 5773 623 5779 717
rect 5821 723 5827 1036
rect 5853 1004 5859 1177
rect 5885 1144 5891 1617
rect 5949 1544 5955 1856
rect 5965 1844 5971 2516
rect 6045 2504 6051 2636
rect 6061 2364 6067 2936
rect 6077 2904 6083 2936
rect 6077 2644 6083 2656
rect 6077 2504 6083 2556
rect 6093 2463 6099 3077
rect 6125 3064 6131 3116
rect 6141 3064 6147 3277
rect 6157 3144 6163 3236
rect 6125 2924 6131 2936
rect 6141 2924 6147 3036
rect 6173 3024 6179 3376
rect 6189 3244 6195 3456
rect 6237 3444 6243 3476
rect 6253 3324 6259 3336
rect 6205 3284 6211 3316
rect 6221 3103 6227 3136
rect 6221 3097 6243 3103
rect 6205 3084 6211 3096
rect 6237 3044 6243 3097
rect 6173 2943 6179 2996
rect 6253 2984 6259 3276
rect 6285 3104 6291 3116
rect 6269 2984 6275 2996
rect 6164 2937 6179 2943
rect 6125 2744 6131 2836
rect 6157 2804 6163 2936
rect 6237 2924 6243 2956
rect 6205 2904 6211 2916
rect 6109 2684 6115 2696
rect 6125 2664 6131 2696
rect 6125 2604 6131 2656
rect 6109 2464 6115 2536
rect 6077 2457 6099 2463
rect 5981 1964 5987 2356
rect 6029 2243 6035 2276
rect 6045 2264 6051 2336
rect 6029 2237 6044 2243
rect 6013 2184 6019 2236
rect 6029 2204 6035 2237
rect 6077 2204 6083 2457
rect 6109 2304 6115 2456
rect 5981 1904 5987 1916
rect 6013 1883 6019 1956
rect 6029 1924 6035 2016
rect 6029 1904 6035 1916
rect 5997 1877 6019 1883
rect 5981 1704 5987 1796
rect 5965 1544 5971 1636
rect 5981 1524 5987 1576
rect 5949 1483 5955 1496
rect 5933 1477 5955 1483
rect 5917 1464 5923 1476
rect 5901 1364 5907 1436
rect 5917 1343 5923 1416
rect 5901 1337 5923 1343
rect 5901 1284 5907 1337
rect 5917 1304 5923 1316
rect 5933 1204 5939 1477
rect 5965 1344 5971 1416
rect 5997 1384 6003 1877
rect 6013 1844 6019 1856
rect 6013 1764 6019 1816
rect 6013 1643 6019 1718
rect 6045 1683 6051 2016
rect 6061 1984 6067 2056
rect 6093 2024 6099 2156
rect 6109 2084 6115 2296
rect 6061 1904 6067 1916
rect 6093 1884 6099 1956
rect 6125 1944 6131 2576
rect 6157 2564 6163 2736
rect 6173 2724 6179 2836
rect 6189 2703 6195 2796
rect 6205 2784 6211 2896
rect 6237 2724 6243 2836
rect 6173 2697 6195 2703
rect 6157 2524 6163 2536
rect 6141 2204 6147 2376
rect 6157 2324 6163 2496
rect 6157 2284 6163 2296
rect 6157 2084 6163 2116
rect 6157 1984 6163 2016
rect 6077 1764 6083 1776
rect 6045 1677 6067 1683
rect 6013 1637 6035 1643
rect 6029 1504 6035 1637
rect 6061 1343 6067 1677
rect 6093 1503 6099 1876
rect 6109 1824 6115 1916
rect 6141 1904 6147 1916
rect 6125 1803 6131 1876
rect 6109 1797 6131 1803
rect 6109 1643 6115 1797
rect 6109 1637 6131 1643
rect 6093 1497 6115 1503
rect 6061 1337 6083 1343
rect 6013 1324 6019 1336
rect 5869 1083 5875 1116
rect 5885 1104 5891 1116
rect 5901 1104 5907 1176
rect 5869 1077 5884 1083
rect 5917 1083 5923 1136
rect 5933 1084 5939 1196
rect 5901 1077 5923 1083
rect 5869 983 5875 1056
rect 5901 983 5907 1077
rect 5853 977 5875 983
rect 5885 977 5907 983
rect 5837 803 5843 876
rect 5853 824 5859 977
rect 5885 884 5891 977
rect 5933 964 5939 1056
rect 5949 984 5955 1236
rect 5981 1223 5987 1276
rect 5997 1244 6003 1316
rect 6029 1304 6035 1316
rect 6077 1303 6083 1337
rect 6061 1297 6083 1303
rect 5981 1217 6003 1223
rect 5965 1064 5971 1176
rect 5997 1103 6003 1217
rect 6013 1184 6019 1196
rect 5981 1097 6003 1103
rect 5981 1084 5987 1097
rect 5965 997 6003 1003
rect 5965 964 5971 997
rect 5997 984 6003 997
rect 5908 957 5923 963
rect 5917 944 5923 957
rect 5981 944 5987 976
rect 5837 797 5875 803
rect 5869 763 5875 797
rect 5885 784 5891 816
rect 5901 764 5907 936
rect 5933 864 5939 916
rect 5965 784 5971 936
rect 5997 924 6003 936
rect 5981 824 5987 916
rect 6013 784 6019 1136
rect 6029 1064 6035 1096
rect 6045 1084 6051 1136
rect 6045 984 6051 1016
rect 6029 884 6035 896
rect 6045 824 6051 956
rect 6061 884 6067 1297
rect 6093 1104 6099 1456
rect 6109 1324 6115 1497
rect 6125 1464 6131 1637
rect 6141 1403 6147 1616
rect 6157 1604 6163 1936
rect 6173 1884 6179 2697
rect 6189 2664 6195 2676
rect 6189 2384 6195 2556
rect 6221 2444 6227 2656
rect 6253 2364 6259 2816
rect 6269 2584 6275 2956
rect 6285 2583 6291 3096
rect 6301 2604 6307 4476
rect 6285 2577 6307 2583
rect 6189 2024 6195 2196
rect 6205 2124 6211 2336
rect 6189 1984 6195 1996
rect 6189 1864 6195 1956
rect 6205 1944 6211 1956
rect 6205 1864 6211 1896
rect 6173 1523 6179 1856
rect 6189 1724 6195 1776
rect 6173 1517 6195 1523
rect 6141 1397 6163 1403
rect 6109 1203 6115 1276
rect 6109 1197 6131 1203
rect 6125 1163 6131 1197
rect 6141 1184 6147 1276
rect 6125 1157 6147 1163
rect 6077 904 6083 1056
rect 6093 1043 6099 1076
rect 6109 1064 6115 1116
rect 6125 1084 6131 1136
rect 6093 1037 6115 1043
rect 6109 964 6115 1037
rect 6077 843 6083 876
rect 6077 837 6099 843
rect 5981 777 6003 783
rect 5869 757 5891 763
rect 5837 724 5843 756
rect 5805 717 5827 723
rect 5773 617 5795 623
rect 5741 583 5747 596
rect 5732 577 5747 583
rect 5725 537 5740 543
rect 5588 517 5603 523
rect 5549 504 5555 516
rect 5565 464 5571 496
rect 5405 284 5411 336
rect 5421 317 5468 323
rect 5421 304 5427 317
rect 5485 304 5491 356
rect 5469 163 5475 296
rect 5501 264 5507 336
rect 5581 324 5587 356
rect 5533 264 5539 316
rect 5597 304 5603 416
rect 5613 304 5619 516
rect 5661 483 5667 536
rect 5725 523 5731 537
rect 5629 477 5667 483
rect 5629 303 5635 477
rect 5645 344 5651 456
rect 5661 443 5667 477
rect 5709 517 5731 523
rect 5709 443 5715 517
rect 5661 437 5715 443
rect 5629 297 5644 303
rect 5485 184 5491 236
rect 5517 164 5523 256
rect 5469 157 5491 163
rect 5453 144 5459 156
rect 5357 137 5379 143
rect 5117 57 5139 63
rect 5133 43 5139 57
rect 5133 37 5276 43
rect 5293 23 5299 116
rect 5309 44 5315 136
rect 5332 117 5340 123
rect 5373 64 5379 137
rect 5469 103 5475 116
rect 5460 97 5475 103
rect 5469 84 5475 97
rect 5485 63 5491 157
rect 5565 104 5571 276
rect 5581 204 5587 296
rect 5645 284 5651 296
rect 5661 263 5667 316
rect 5677 284 5683 376
rect 5693 303 5699 396
rect 5709 324 5715 396
rect 5725 384 5731 496
rect 5725 304 5731 336
rect 5693 297 5715 303
rect 5709 284 5715 297
rect 5725 263 5731 276
rect 5629 257 5667 263
rect 5677 257 5731 263
rect 5629 104 5635 257
rect 5677 243 5683 257
rect 5652 237 5683 243
rect 5693 203 5699 236
rect 5677 197 5699 203
rect 5661 124 5667 176
rect 5581 83 5587 96
rect 5556 77 5587 83
rect 5677 64 5683 197
rect 5741 184 5747 476
rect 5773 383 5779 576
rect 5789 524 5795 617
rect 5805 584 5811 717
rect 5869 723 5875 736
rect 5853 717 5875 723
rect 5853 704 5859 717
rect 5844 677 5875 683
rect 5869 604 5875 677
rect 5885 664 5891 757
rect 5917 684 5923 776
rect 5805 544 5811 556
rect 5789 484 5795 516
rect 5757 377 5779 383
rect 5757 184 5763 377
rect 5789 344 5795 356
rect 5773 264 5779 316
rect 5789 304 5795 336
rect 5469 57 5491 63
rect 5357 23 5363 36
rect 5469 24 5475 57
rect 5757 24 5763 156
rect 5789 44 5795 276
rect 5837 204 5843 596
rect 5885 584 5891 596
rect 5901 564 5907 676
rect 5917 564 5923 636
rect 5933 604 5939 776
rect 5981 763 5987 777
rect 5965 757 5987 763
rect 5997 763 6003 777
rect 5997 757 6019 763
rect 5965 703 5971 757
rect 6013 704 6019 757
rect 6077 704 6083 796
rect 6093 784 6099 837
rect 5956 697 5971 703
rect 5997 664 6003 676
rect 6093 664 6099 756
rect 6109 724 6115 896
rect 6125 683 6131 1056
rect 6141 944 6147 1157
rect 6109 677 6131 683
rect 5933 564 5939 596
rect 5949 584 5955 656
rect 5965 544 5971 656
rect 5853 524 5859 536
rect 5869 524 5875 536
rect 5917 504 5923 516
rect 5997 504 6003 596
rect 6077 584 6083 656
rect 6077 564 6083 576
rect 6061 523 6067 556
rect 6061 517 6076 523
rect 5853 364 5859 436
rect 5853 324 5859 336
rect 5885 264 5891 316
rect 5933 304 5939 336
rect 5965 284 5971 496
rect 5853 84 5859 256
rect 5901 243 5907 256
rect 5885 237 5907 243
rect 5885 104 5891 237
rect 5965 184 5971 236
rect 5981 124 5987 396
rect 6013 364 6019 496
rect 6013 304 6019 336
rect 6029 304 6035 396
rect 6061 324 6067 336
rect 5997 184 6003 276
rect 6029 264 6035 296
rect 6045 264 6051 276
rect 6045 224 6051 256
rect 6061 204 6067 296
rect 6077 224 6083 456
rect 6093 444 6099 656
rect 6109 624 6115 677
rect 6125 584 6131 636
rect 6141 584 6147 936
rect 6157 744 6163 1397
rect 6173 1184 6179 1476
rect 6189 1384 6195 1517
rect 6205 1504 6211 1816
rect 6221 1804 6227 2236
rect 6237 2203 6243 2256
rect 6253 2224 6259 2296
rect 6237 2197 6259 2203
rect 6253 1924 6259 2197
rect 6269 2184 6275 2476
rect 6269 1964 6275 2076
rect 6301 2004 6307 2577
rect 6253 1884 6259 1896
rect 6221 1504 6227 1536
rect 6205 1424 6211 1476
rect 6205 1364 6211 1416
rect 6189 1304 6195 1316
rect 6189 1204 6195 1276
rect 6205 1124 6211 1196
rect 6189 1084 6195 1116
rect 6173 926 6179 976
rect 6237 964 6243 1876
rect 6269 1284 6275 1596
rect 6269 1103 6275 1256
rect 6253 1097 6275 1103
rect 6253 964 6259 1097
rect 6173 917 6179 918
rect 6205 723 6211 956
rect 6237 744 6243 836
rect 6253 764 6259 876
rect 6189 717 6211 723
rect 6157 704 6163 716
rect 6173 683 6179 716
rect 6157 677 6179 683
rect 6157 564 6163 677
rect 6093 324 6099 356
rect 6093 284 6099 316
rect 6109 304 6115 396
rect 6141 384 6147 476
rect 6189 383 6195 717
rect 6253 704 6259 716
rect 6205 584 6211 676
rect 6205 484 6211 556
rect 6221 424 6227 616
rect 6253 584 6259 676
rect 6253 544 6259 576
rect 6269 504 6275 1016
rect 6285 924 6291 1076
rect 6285 877 6300 883
rect 6285 844 6291 877
rect 6285 784 6291 816
rect 6285 564 6291 736
rect 6189 377 6211 383
rect 6141 324 6147 376
rect 6109 264 6115 276
rect 6125 264 6131 276
rect 6109 144 6115 256
rect 6157 244 6163 316
rect 6157 184 6163 216
rect 6189 184 6195 356
rect 6205 204 6211 377
rect 6173 164 6179 176
rect 6260 157 6268 163
rect 6221 144 6227 156
rect 5901 104 5907 118
rect 6029 64 6035 116
rect 5293 17 5363 23
rect 4637 -23 4739 -17
rect 3245 -43 3299 -37
<< m3contact >>
rect 396 4596 404 4604
rect 44 4536 52 4544
rect 108 4536 116 4544
rect 12 4516 20 4524
rect 92 4516 100 4524
rect 252 4516 260 4524
rect 12 4356 20 4364
rect 140 4302 148 4304
rect 140 4296 148 4302
rect 172 4296 180 4304
rect 124 4136 132 4144
rect 76 4056 84 4064
rect 476 4516 484 4524
rect 364 4456 372 4464
rect 460 4456 468 4464
rect 204 4196 212 4204
rect 188 4176 196 4184
rect 668 4576 676 4584
rect 732 4576 740 4584
rect 668 4516 676 4524
rect 620 4496 628 4504
rect 716 4496 724 4504
rect 732 4456 740 4464
rect 620 4296 628 4304
rect 396 4196 404 4204
rect 380 4176 388 4184
rect 284 4156 292 4164
rect 332 4156 340 4164
rect 188 4116 196 4124
rect 204 4076 212 4084
rect 332 4096 340 4104
rect 348 4096 356 4104
rect 572 4176 580 4184
rect 652 4176 660 4184
rect 428 4156 436 4164
rect 476 4156 484 4164
rect 700 4156 708 4164
rect 556 4136 564 4144
rect 668 4136 676 4144
rect 412 4116 420 4124
rect 396 4096 404 4104
rect 316 4076 324 4084
rect 364 4076 372 4084
rect 364 4056 372 4064
rect 748 4116 756 4124
rect 604 4096 612 4104
rect 636 4096 644 4104
rect 76 3956 84 3964
rect 268 3956 276 3964
rect 284 3956 292 3964
rect 252 3936 260 3944
rect 92 3916 100 3924
rect 332 3936 340 3944
rect 76 3896 84 3904
rect 124 3896 132 3904
rect 284 3896 292 3904
rect 108 3876 116 3884
rect 412 3916 420 3924
rect 524 3916 532 3924
rect 348 3896 356 3904
rect 156 3876 164 3884
rect 172 3876 180 3884
rect 204 3876 212 3884
rect 252 3876 260 3884
rect 156 3856 164 3864
rect 140 3836 148 3844
rect 220 3856 228 3864
rect 236 3836 244 3844
rect 316 3836 324 3844
rect 252 3816 260 3824
rect 236 3796 244 3804
rect 44 3776 52 3784
rect 92 3776 100 3784
rect 124 3776 132 3784
rect 204 3776 212 3784
rect 332 3796 340 3804
rect 284 3776 292 3784
rect 300 3776 308 3784
rect 60 3736 68 3744
rect 92 3736 100 3744
rect 124 3736 132 3744
rect 28 3636 36 3644
rect 76 3716 84 3724
rect 92 3716 100 3724
rect 124 3716 132 3724
rect 140 3716 148 3724
rect 140 3696 148 3704
rect 44 3596 52 3604
rect 76 3596 84 3604
rect 124 3596 132 3604
rect 316 3736 324 3744
rect 268 3716 276 3724
rect 300 3656 308 3664
rect 332 3636 340 3644
rect 204 3596 212 3604
rect 412 3896 420 3904
rect 364 3836 372 3844
rect 380 3836 388 3844
rect 460 3876 468 3884
rect 508 3856 516 3864
rect 508 3836 516 3844
rect 460 3796 468 3804
rect 364 3736 372 3744
rect 396 3716 404 3724
rect 412 3716 420 3724
rect 476 3736 484 3744
rect 492 3736 500 3744
rect 860 4516 868 4524
rect 844 4456 852 4464
rect 1020 4576 1028 4584
rect 972 4556 980 4564
rect 1068 4576 1076 4584
rect 1100 4516 1108 4524
rect 1020 4496 1028 4504
rect 1084 4496 1092 4504
rect 1036 4476 1044 4484
rect 1116 4476 1124 4484
rect 1084 4436 1092 4444
rect 940 4336 948 4344
rect 1036 4336 1044 4344
rect 1260 4556 1268 4564
rect 1372 4536 1380 4544
rect 1340 4476 1348 4484
rect 1244 4456 1252 4464
rect 1276 4456 1284 4464
rect 828 4296 836 4304
rect 1004 4296 1012 4304
rect 1036 4296 1044 4304
rect 1084 4296 1092 4304
rect 1196 4296 1204 4304
rect 812 4216 820 4224
rect 876 4256 884 4264
rect 860 4196 868 4204
rect 892 4156 900 4164
rect 908 4136 916 4144
rect 876 4076 884 4084
rect 988 4256 996 4264
rect 1068 4256 1076 4264
rect 1116 4256 1124 4264
rect 956 4176 964 4184
rect 972 4156 980 4164
rect 956 4136 964 4144
rect 1052 4196 1060 4204
rect 1020 4136 1028 4144
rect 1100 4216 1108 4224
rect 1100 4156 1108 4164
rect 988 4116 996 4124
rect 1004 4116 1012 4124
rect 1036 4116 1044 4124
rect 1084 4116 1092 4124
rect 924 4076 932 4084
rect 988 4096 996 4104
rect 988 4076 996 4084
rect 908 4056 916 4064
rect 972 4056 980 4064
rect 876 4016 884 4024
rect 780 3996 788 4004
rect 684 3916 692 3924
rect 572 3876 580 3884
rect 636 3876 644 3884
rect 588 3776 596 3784
rect 524 3756 532 3764
rect 540 3736 548 3744
rect 540 3716 548 3724
rect 524 3696 532 3704
rect 540 3696 548 3704
rect 588 3696 596 3704
rect 396 3676 404 3684
rect 428 3636 436 3644
rect 76 3556 84 3564
rect 204 3556 212 3564
rect 348 3556 356 3564
rect 284 3536 292 3544
rect 60 3516 68 3524
rect 44 3496 52 3504
rect 76 3496 84 3504
rect 124 3496 132 3504
rect 172 3496 180 3504
rect 44 3476 52 3484
rect 188 3476 196 3484
rect 140 3456 148 3464
rect 220 3476 228 3484
rect 412 3516 420 3524
rect 316 3496 324 3504
rect 396 3496 404 3504
rect 492 3596 500 3604
rect 348 3476 356 3484
rect 396 3476 404 3484
rect 428 3476 436 3484
rect 492 3476 500 3484
rect 220 3456 228 3464
rect 172 3436 180 3444
rect 204 3436 212 3444
rect 124 3376 132 3384
rect 188 3356 196 3364
rect 172 3316 180 3324
rect 188 3176 196 3184
rect 332 3396 340 3404
rect 556 3676 564 3684
rect 860 3916 868 3924
rect 860 3896 868 3904
rect 844 3876 852 3884
rect 636 3816 644 3824
rect 700 3796 708 3804
rect 812 3796 820 3804
rect 844 3776 852 3784
rect 892 3936 900 3944
rect 828 3736 836 3744
rect 860 3736 868 3744
rect 812 3716 820 3724
rect 636 3696 644 3704
rect 668 3696 676 3704
rect 572 3576 580 3584
rect 556 3516 564 3524
rect 572 3516 580 3524
rect 540 3476 548 3484
rect 572 3476 580 3484
rect 572 3456 580 3464
rect 364 3376 372 3384
rect 428 3336 436 3344
rect 268 3316 276 3324
rect 300 3318 308 3324
rect 300 3316 308 3318
rect 540 3396 548 3404
rect 508 3356 516 3364
rect 556 3356 564 3364
rect 556 3336 564 3344
rect 476 3316 484 3324
rect 220 3256 228 3264
rect 204 3156 212 3164
rect 92 3116 100 3124
rect 220 3116 228 3124
rect 220 3096 228 3104
rect 204 3056 212 3064
rect 460 3276 468 3284
rect 348 3216 356 3224
rect 444 3216 452 3224
rect 412 3196 420 3204
rect 364 3156 372 3164
rect 412 3156 420 3164
rect 316 3136 324 3144
rect 428 3136 436 3144
rect 460 3136 468 3144
rect 348 3116 356 3124
rect 252 3096 260 3104
rect 284 3096 292 3104
rect 284 3036 292 3044
rect 300 3036 308 3044
rect 236 2976 244 2984
rect 28 2956 36 2964
rect 60 2916 68 2924
rect 12 2896 20 2904
rect 76 2856 84 2864
rect 156 2916 164 2924
rect 156 2896 164 2904
rect 348 2976 356 2984
rect 332 2936 340 2944
rect 380 2936 388 2944
rect 220 2896 228 2904
rect 284 2876 292 2884
rect 140 2856 148 2864
rect 188 2856 196 2864
rect 252 2856 260 2864
rect 316 2836 324 2844
rect 492 3296 500 3304
rect 524 3256 532 3264
rect 492 3116 500 3124
rect 540 3196 548 3204
rect 524 3096 532 3104
rect 508 3016 516 3024
rect 508 2936 516 2944
rect 492 2916 500 2924
rect 364 2896 372 2904
rect 396 2896 404 2904
rect 412 2896 420 2904
rect 396 2856 404 2864
rect 124 2776 132 2784
rect 140 2776 148 2784
rect 220 2776 228 2784
rect 92 2736 100 2744
rect 76 2696 84 2704
rect 220 2756 228 2764
rect 236 2756 244 2764
rect 156 2716 164 2724
rect 188 2716 196 2724
rect 172 2696 180 2704
rect 252 2736 260 2744
rect 268 2696 276 2704
rect 172 2676 180 2684
rect 220 2676 228 2684
rect 92 2576 100 2584
rect 44 2556 52 2564
rect 12 2536 20 2544
rect 44 2536 52 2544
rect 92 2536 100 2544
rect 140 2536 148 2544
rect 28 2516 36 2524
rect 124 2516 132 2524
rect 252 2616 260 2624
rect 284 2616 292 2624
rect 332 2716 340 2724
rect 364 2696 372 2704
rect 300 2596 308 2604
rect 620 3636 628 3644
rect 604 3616 612 3624
rect 652 3596 660 3604
rect 636 3576 644 3584
rect 604 3516 612 3524
rect 604 3496 612 3504
rect 636 3496 644 3504
rect 748 3596 756 3604
rect 764 3596 772 3604
rect 700 3516 708 3524
rect 684 3496 692 3504
rect 604 3476 612 3484
rect 588 3336 596 3344
rect 620 3456 628 3464
rect 652 3456 660 3464
rect 764 3536 772 3544
rect 796 3536 804 3544
rect 876 3716 884 3724
rect 876 3596 884 3604
rect 988 4036 996 4044
rect 940 3996 948 4004
rect 908 3896 916 3904
rect 1020 4076 1028 4084
rect 1100 4076 1108 4084
rect 1084 4056 1092 4064
rect 1148 4056 1156 4064
rect 1116 4036 1124 4044
rect 1036 3976 1044 3984
rect 1116 3976 1124 3984
rect 1132 3976 1140 3984
rect 1020 3916 1028 3924
rect 1004 3896 1012 3904
rect 956 3856 964 3864
rect 908 3836 916 3844
rect 924 3736 932 3744
rect 956 3736 964 3744
rect 908 3696 916 3704
rect 940 3676 948 3684
rect 908 3656 916 3664
rect 1004 3716 1012 3724
rect 988 3676 996 3684
rect 972 3656 980 3664
rect 956 3556 964 3564
rect 860 3536 868 3544
rect 892 3536 900 3544
rect 812 3496 820 3504
rect 780 3476 788 3484
rect 796 3476 804 3484
rect 620 3396 628 3404
rect 684 3376 692 3384
rect 668 3356 676 3364
rect 636 3336 644 3344
rect 780 3336 788 3344
rect 604 3316 612 3324
rect 636 3316 644 3324
rect 684 3316 692 3324
rect 716 3316 724 3324
rect 764 3316 772 3324
rect 588 3296 596 3304
rect 668 3296 676 3304
rect 716 3296 724 3304
rect 748 3296 756 3304
rect 588 3276 596 3284
rect 604 3236 612 3244
rect 684 3236 692 3244
rect 716 3236 724 3244
rect 588 3196 596 3204
rect 588 3176 596 3184
rect 604 3156 612 3164
rect 556 3116 564 3124
rect 572 3116 580 3124
rect 572 3096 580 3104
rect 652 3116 660 3124
rect 732 3156 740 3164
rect 716 3136 724 3144
rect 716 3116 724 3124
rect 572 3076 580 3084
rect 620 3076 628 3084
rect 684 3076 692 3084
rect 556 3056 564 3064
rect 540 2996 548 3004
rect 540 2956 548 2964
rect 556 2936 564 2944
rect 540 2916 548 2924
rect 524 2836 532 2844
rect 412 2756 420 2764
rect 428 2736 436 2744
rect 444 2736 452 2744
rect 412 2696 420 2704
rect 460 2696 468 2704
rect 524 2756 532 2764
rect 700 3056 708 3064
rect 636 3036 644 3044
rect 620 3016 628 3024
rect 604 2956 612 2964
rect 572 2916 580 2924
rect 588 2856 596 2864
rect 604 2836 612 2844
rect 572 2796 580 2804
rect 556 2756 564 2764
rect 540 2716 548 2724
rect 588 2716 596 2724
rect 380 2676 388 2684
rect 428 2636 436 2644
rect 348 2596 356 2604
rect 316 2576 324 2584
rect 332 2576 340 2584
rect 364 2536 372 2544
rect 284 2516 292 2524
rect 300 2516 308 2524
rect 140 2376 148 2384
rect 348 2336 356 2344
rect 300 2316 308 2324
rect 332 2316 340 2324
rect 12 2296 20 2304
rect 188 2296 196 2304
rect 60 2276 68 2284
rect 300 2276 308 2284
rect 140 2256 148 2264
rect 332 2256 340 2264
rect 444 2616 452 2624
rect 396 2518 404 2524
rect 396 2516 404 2518
rect 428 2516 436 2524
rect 412 2356 420 2364
rect 380 2276 388 2284
rect 428 2316 436 2324
rect 508 2676 516 2684
rect 492 2636 500 2644
rect 508 2616 516 2624
rect 508 2576 516 2584
rect 460 2556 468 2564
rect 492 2556 500 2564
rect 460 2536 468 2544
rect 476 2396 484 2404
rect 508 2356 516 2364
rect 428 2236 436 2244
rect 396 2216 404 2224
rect 364 2196 372 2204
rect 140 2156 148 2164
rect 204 2156 212 2164
rect 252 2156 260 2164
rect 300 2156 308 2164
rect 348 2156 356 2164
rect 428 2156 436 2164
rect 124 2136 132 2144
rect 76 2096 84 2104
rect 12 1996 20 2004
rect 108 1896 116 1904
rect 60 1756 68 1764
rect 28 1736 36 1744
rect 316 2116 324 2124
rect 204 2096 212 2104
rect 140 1916 148 1924
rect 204 1896 212 1904
rect 236 1896 244 1904
rect 172 1876 180 1884
rect 172 1856 180 1864
rect 220 1856 228 1864
rect 188 1836 196 1844
rect 124 1736 132 1744
rect 172 1736 180 1744
rect 12 1716 20 1724
rect 108 1716 116 1724
rect 252 1836 260 1844
rect 236 1756 244 1764
rect 108 1696 116 1704
rect 156 1696 164 1704
rect 172 1696 180 1704
rect 204 1696 212 1704
rect 44 1496 52 1504
rect 220 1496 228 1504
rect 204 1476 212 1484
rect 572 2656 580 2664
rect 652 2956 660 2964
rect 780 3156 788 3164
rect 892 3516 900 3524
rect 844 3476 852 3484
rect 860 3476 868 3484
rect 892 3476 900 3484
rect 828 3456 836 3464
rect 828 3356 836 3364
rect 828 3316 836 3324
rect 844 3316 852 3324
rect 844 3296 852 3304
rect 1068 3956 1076 3964
rect 1084 3896 1092 3904
rect 1068 3876 1076 3884
rect 1084 3876 1092 3884
rect 1084 3856 1092 3864
rect 1148 3916 1156 3924
rect 1276 4276 1284 4284
rect 1260 4216 1268 4224
rect 1244 4116 1252 4124
rect 1292 4236 1300 4244
rect 1324 4236 1332 4244
rect 1548 4616 1556 4624
rect 1628 4616 1636 4624
rect 1708 4616 1716 4624
rect 1724 4616 1732 4624
rect 1756 4616 1764 4624
rect 1420 4496 1428 4504
rect 1516 4518 1524 4524
rect 1516 4516 1524 4518
rect 1500 4456 1508 4464
rect 1580 4536 1588 4544
rect 1596 4536 1604 4544
rect 1788 4536 1796 4544
rect 1596 4496 1604 4504
rect 1644 4516 1652 4524
rect 1676 4516 1684 4524
rect 1628 4496 1636 4504
rect 1660 4476 1668 4484
rect 1676 4476 1684 4484
rect 1612 4436 1620 4444
rect 1644 4436 1652 4444
rect 1577 4406 1585 4414
rect 1587 4406 1595 4414
rect 1597 4406 1605 4414
rect 1607 4406 1615 4414
rect 1532 4376 1540 4384
rect 1548 4376 1556 4384
rect 1580 4376 1588 4384
rect 1484 4336 1492 4344
rect 1372 4276 1380 4284
rect 1356 4236 1364 4244
rect 1532 4316 1540 4324
rect 1452 4276 1460 4284
rect 1500 4276 1508 4284
rect 1404 4256 1412 4264
rect 1484 4256 1492 4264
rect 1532 4256 1540 4264
rect 1468 4216 1476 4224
rect 1436 4136 1444 4144
rect 1340 4116 1348 4124
rect 1308 4096 1316 4104
rect 1356 4096 1364 4104
rect 1212 4056 1220 4064
rect 1356 4056 1364 4064
rect 1388 4056 1396 4064
rect 1196 4016 1204 4024
rect 1340 4016 1348 4024
rect 1292 3996 1300 4004
rect 1180 3976 1188 3984
rect 1180 3916 1188 3924
rect 1228 3916 1236 3924
rect 1244 3916 1252 3924
rect 1132 3856 1140 3864
rect 1116 3776 1124 3784
rect 1084 3756 1092 3764
rect 1100 3756 1108 3764
rect 1068 3736 1076 3744
rect 1260 3856 1268 3864
rect 1468 4096 1476 4104
rect 1692 4416 1700 4424
rect 1660 4356 1668 4364
rect 1548 4216 1556 4224
rect 1500 4136 1508 4144
rect 1452 4016 1460 4024
rect 1388 3996 1396 4004
rect 1436 3996 1444 4004
rect 1452 3996 1460 4004
rect 1404 3936 1412 3944
rect 1356 3876 1364 3884
rect 1436 3876 1444 3884
rect 1164 3836 1172 3844
rect 1196 3836 1204 3844
rect 1116 3736 1124 3744
rect 1132 3736 1140 3744
rect 1148 3736 1156 3744
rect 1276 3776 1284 3784
rect 1052 3696 1060 3704
rect 1068 3696 1076 3704
rect 1036 3636 1044 3644
rect 1036 3616 1044 3624
rect 1052 3616 1060 3624
rect 1004 3536 1012 3544
rect 972 3516 980 3524
rect 972 3476 980 3484
rect 1052 3556 1060 3564
rect 1116 3696 1124 3704
rect 1100 3676 1108 3684
rect 1084 3596 1092 3604
rect 1084 3576 1092 3584
rect 1020 3476 1028 3484
rect 1148 3716 1156 3724
rect 1228 3716 1236 3724
rect 1132 3576 1140 3584
rect 1116 3556 1124 3564
rect 1116 3536 1124 3544
rect 1340 3836 1348 3844
rect 1436 3836 1444 3844
rect 1452 3836 1460 3844
rect 1580 4256 1588 4264
rect 1596 4256 1604 4264
rect 1740 4516 1748 4524
rect 1740 4496 1748 4504
rect 1788 4496 1796 4504
rect 1756 4356 1764 4364
rect 1772 4356 1780 4364
rect 1628 4176 1636 4184
rect 1692 4176 1700 4184
rect 1788 4316 1796 4324
rect 1596 4156 1604 4164
rect 1612 4156 1620 4164
rect 1548 4096 1556 4104
rect 1532 4056 1540 4064
rect 1548 4056 1556 4064
rect 1516 4016 1524 4024
rect 1676 4156 1684 4164
rect 1740 4156 1748 4164
rect 1644 4096 1652 4104
rect 1577 4006 1585 4014
rect 1587 4006 1595 4014
rect 1597 4006 1605 4014
rect 1607 4006 1615 4014
rect 1596 3896 1604 3904
rect 1484 3856 1492 3864
rect 1500 3816 1508 3824
rect 1436 3756 1444 3764
rect 1468 3756 1476 3764
rect 1372 3736 1380 3744
rect 1388 3736 1396 3744
rect 1244 3696 1252 3704
rect 1260 3696 1268 3704
rect 1164 3676 1172 3684
rect 1180 3676 1188 3684
rect 1180 3616 1188 3624
rect 1212 3576 1220 3584
rect 1180 3556 1188 3564
rect 1196 3556 1204 3564
rect 1116 3516 1124 3524
rect 1148 3516 1156 3524
rect 1180 3516 1188 3524
rect 1100 3476 1108 3484
rect 1020 3456 1028 3464
rect 924 3416 932 3424
rect 956 3396 964 3404
rect 892 3376 900 3384
rect 908 3376 916 3384
rect 940 3376 948 3384
rect 1004 3416 1012 3424
rect 1036 3416 1044 3424
rect 908 3316 916 3324
rect 972 3316 980 3324
rect 988 3316 996 3324
rect 972 3296 980 3304
rect 876 3256 884 3264
rect 876 3236 884 3244
rect 844 3196 852 3204
rect 876 3196 884 3204
rect 748 3076 756 3084
rect 764 3056 772 3064
rect 812 3096 820 3104
rect 700 2956 708 2964
rect 732 2956 740 2964
rect 796 2956 804 2964
rect 812 2956 820 2964
rect 1196 3476 1204 3484
rect 1228 3536 1236 3544
rect 1244 3516 1252 3524
rect 1308 3536 1316 3544
rect 1292 3516 1300 3524
rect 1260 3496 1268 3504
rect 1276 3496 1284 3504
rect 1292 3476 1300 3484
rect 1100 3456 1108 3464
rect 1132 3456 1140 3464
rect 1180 3456 1188 3464
rect 1020 3396 1028 3404
rect 1068 3396 1076 3404
rect 1100 3396 1108 3404
rect 1116 3396 1124 3404
rect 1004 3136 1012 3144
rect 908 3116 916 3124
rect 940 3116 948 3124
rect 988 3116 996 3124
rect 860 3076 868 3084
rect 908 3076 916 3084
rect 748 2916 756 2924
rect 844 2916 852 2924
rect 732 2896 736 2904
rect 736 2896 740 2904
rect 716 2876 724 2884
rect 668 2776 676 2784
rect 668 2756 676 2764
rect 636 2716 644 2724
rect 748 2716 756 2724
rect 716 2676 724 2684
rect 652 2656 660 2664
rect 620 2616 628 2624
rect 684 2616 692 2624
rect 604 2576 612 2584
rect 556 2556 564 2564
rect 540 2516 548 2524
rect 540 2496 548 2504
rect 540 2476 548 2484
rect 524 2336 532 2344
rect 524 2316 532 2324
rect 540 2316 548 2324
rect 572 2536 580 2544
rect 572 2516 580 2524
rect 588 2496 596 2504
rect 572 2296 580 2304
rect 540 2276 548 2284
rect 556 2276 564 2284
rect 524 2236 532 2244
rect 300 2096 308 2104
rect 396 2116 404 2124
rect 460 2116 468 2124
rect 524 2136 532 2144
rect 572 2256 580 2264
rect 428 2056 436 2064
rect 396 2016 404 2024
rect 348 1976 356 1984
rect 284 1916 292 1924
rect 412 1996 420 2004
rect 428 1956 436 1964
rect 444 1936 452 1944
rect 428 1916 436 1924
rect 284 1896 292 1904
rect 380 1896 388 1904
rect 364 1876 372 1884
rect 332 1756 340 1764
rect 556 2096 564 2104
rect 572 2096 580 2104
rect 476 2076 484 2084
rect 620 2556 628 2564
rect 748 2556 756 2564
rect 732 2516 740 2524
rect 652 2496 660 2504
rect 652 2456 660 2464
rect 636 2396 644 2404
rect 620 2356 628 2364
rect 716 2496 724 2504
rect 684 2476 692 2484
rect 668 2416 676 2424
rect 668 2356 676 2364
rect 652 2336 660 2344
rect 636 2296 644 2304
rect 780 2496 788 2504
rect 764 2436 772 2444
rect 764 2416 772 2424
rect 796 2396 804 2404
rect 764 2376 772 2384
rect 748 2356 756 2364
rect 732 2316 740 2324
rect 652 2276 660 2284
rect 684 2276 692 2284
rect 620 2256 628 2264
rect 684 2216 692 2224
rect 1036 3376 1044 3384
rect 1068 3356 1076 3364
rect 1052 3316 1060 3324
rect 1084 3316 1092 3324
rect 988 3096 996 3104
rect 1020 3096 1028 3104
rect 876 3056 884 3064
rect 924 3056 932 3064
rect 956 3056 964 3064
rect 876 3016 884 3024
rect 924 3016 932 3024
rect 940 3016 948 3024
rect 876 2896 884 2904
rect 1020 3076 1028 3084
rect 972 3016 980 3024
rect 1004 3016 1012 3024
rect 956 2896 964 2904
rect 956 2876 964 2884
rect 908 2856 916 2864
rect 988 2896 996 2904
rect 1180 3396 1188 3404
rect 1164 3356 1172 3364
rect 1260 3396 1268 3404
rect 1244 3376 1252 3384
rect 1276 3376 1284 3384
rect 1340 3596 1348 3604
rect 1356 3556 1364 3564
rect 1340 3516 1348 3524
rect 1404 3696 1412 3704
rect 1372 3536 1380 3544
rect 1468 3736 1476 3744
rect 1484 3736 1492 3744
rect 1468 3716 1476 3724
rect 1484 3716 1492 3724
rect 1452 3676 1460 3684
rect 1484 3676 1492 3684
rect 1468 3596 1476 3604
rect 1436 3556 1444 3564
rect 1420 3516 1428 3524
rect 1404 3496 1412 3504
rect 1372 3476 1380 3484
rect 1436 3476 1444 3484
rect 1356 3456 1364 3464
rect 1372 3456 1380 3464
rect 1324 3416 1332 3424
rect 1116 3316 1124 3324
rect 1068 3276 1076 3284
rect 1100 3276 1108 3284
rect 1084 3236 1092 3244
rect 1132 3236 1140 3244
rect 1116 3196 1124 3204
rect 1068 3176 1076 3184
rect 1068 3116 1076 3124
rect 1164 3296 1172 3304
rect 1180 3296 1188 3304
rect 1148 3176 1156 3184
rect 1308 3356 1316 3364
rect 1244 3336 1252 3344
rect 1276 3316 1284 3324
rect 1292 3296 1300 3304
rect 1196 3216 1204 3224
rect 1244 3196 1252 3204
rect 1196 3156 1204 3164
rect 1148 3116 1156 3124
rect 1180 3116 1188 3124
rect 1164 3096 1172 3104
rect 1196 3096 1204 3104
rect 1228 3156 1236 3164
rect 1308 3176 1316 3184
rect 1356 3296 1364 3304
rect 1436 3396 1444 3404
rect 1420 3316 1428 3324
rect 1404 3276 1412 3284
rect 1356 3256 1364 3264
rect 1388 3256 1396 3264
rect 1356 3216 1364 3224
rect 1244 3136 1252 3144
rect 1228 3116 1236 3124
rect 1260 3116 1268 3124
rect 1148 3076 1156 3084
rect 1132 3036 1140 3044
rect 1084 3016 1092 3024
rect 1116 3016 1124 3024
rect 1052 2956 1060 2964
rect 1036 2936 1044 2944
rect 1116 2936 1124 2944
rect 1020 2916 1028 2924
rect 1084 2916 1092 2924
rect 1148 2956 1156 2964
rect 1036 2896 1044 2904
rect 1100 2896 1108 2904
rect 1132 2896 1140 2904
rect 972 2856 980 2864
rect 1132 2856 1140 2864
rect 892 2816 900 2824
rect 924 2816 932 2824
rect 956 2816 964 2824
rect 892 2776 900 2784
rect 892 2756 900 2764
rect 876 2716 884 2724
rect 908 2716 916 2724
rect 860 2676 868 2684
rect 1100 2836 1108 2844
rect 972 2796 980 2804
rect 1068 2796 1076 2804
rect 940 2736 948 2744
rect 956 2736 964 2744
rect 1116 2816 1124 2824
rect 1116 2736 1124 2744
rect 956 2716 964 2724
rect 1196 3076 1204 3084
rect 1212 3076 1220 3084
rect 1180 3036 1188 3044
rect 1180 2876 1188 2884
rect 1164 2836 1172 2844
rect 1148 2816 1156 2824
rect 1148 2736 1156 2744
rect 956 2696 964 2704
rect 1004 2696 1012 2704
rect 1052 2696 1060 2704
rect 1084 2696 1092 2704
rect 1100 2696 1108 2704
rect 1052 2676 1060 2684
rect 1068 2676 1076 2684
rect 924 2616 932 2624
rect 988 2596 996 2604
rect 940 2556 948 2564
rect 844 2536 852 2544
rect 876 2536 884 2544
rect 972 2536 980 2544
rect 988 2536 996 2544
rect 828 2416 836 2424
rect 876 2496 884 2504
rect 876 2456 884 2464
rect 892 2456 900 2464
rect 1020 2496 1028 2504
rect 988 2476 996 2484
rect 908 2416 916 2424
rect 940 2416 948 2424
rect 812 2376 820 2384
rect 828 2356 836 2364
rect 924 2356 932 2364
rect 844 2316 852 2324
rect 860 2316 868 2324
rect 892 2316 900 2324
rect 892 2296 900 2304
rect 908 2296 916 2304
rect 780 2276 788 2284
rect 940 2336 948 2344
rect 956 2296 964 2304
rect 972 2296 980 2304
rect 940 2276 948 2284
rect 1180 2816 1188 2824
rect 1180 2736 1188 2744
rect 1212 2976 1220 2984
rect 1244 3096 1252 3104
rect 1276 3096 1284 3104
rect 1308 3056 1316 3064
rect 1388 3096 1396 3104
rect 1356 3036 1364 3044
rect 1212 2936 1220 2944
rect 1308 2936 1316 2944
rect 1388 3016 1396 3024
rect 1388 2956 1396 2964
rect 1372 2936 1380 2944
rect 1244 2916 1252 2924
rect 1340 2896 1348 2904
rect 1212 2756 1220 2764
rect 1228 2716 1236 2724
rect 1132 2616 1140 2624
rect 1100 2576 1108 2584
rect 1116 2576 1124 2584
rect 1244 2676 1252 2684
rect 1324 2796 1332 2804
rect 1308 2776 1316 2784
rect 1324 2756 1332 2764
rect 1292 2676 1300 2684
rect 1228 2656 1236 2664
rect 1244 2656 1252 2664
rect 1276 2656 1284 2664
rect 1292 2656 1300 2664
rect 1180 2576 1188 2584
rect 1164 2516 1172 2524
rect 1100 2496 1108 2504
rect 1148 2496 1156 2504
rect 1068 2476 1076 2484
rect 1036 2316 1044 2324
rect 796 2236 804 2244
rect 1020 2256 1028 2264
rect 796 2216 804 2224
rect 812 2216 820 2224
rect 812 2196 820 2204
rect 812 2156 820 2164
rect 716 2096 724 2104
rect 732 2096 740 2104
rect 492 2056 500 2064
rect 556 2056 564 2064
rect 604 2056 612 2064
rect 764 2056 772 2064
rect 476 2016 484 2024
rect 492 2016 500 2024
rect 508 2016 516 2024
rect 476 1996 484 2004
rect 492 1976 500 1984
rect 540 1976 548 1984
rect 396 1836 404 1844
rect 476 1796 484 1804
rect 428 1776 436 1784
rect 780 2016 788 2024
rect 620 1976 628 1984
rect 636 1976 644 1984
rect 668 1976 676 1984
rect 572 1936 580 1944
rect 588 1916 596 1924
rect 476 1756 484 1764
rect 508 1756 516 1764
rect 460 1736 468 1744
rect 316 1716 324 1724
rect 492 1716 500 1724
rect 556 1816 564 1824
rect 300 1636 308 1644
rect 268 1536 276 1544
rect 428 1696 436 1704
rect 524 1616 532 1624
rect 316 1556 324 1564
rect 364 1536 372 1544
rect 300 1516 308 1524
rect 268 1476 276 1484
rect 332 1476 340 1484
rect 316 1416 324 1424
rect 60 1376 68 1384
rect 236 1376 244 1384
rect 156 1356 164 1364
rect 332 1356 340 1364
rect 188 1336 196 1344
rect 316 1336 324 1344
rect 12 1316 20 1324
rect 220 1316 228 1324
rect 156 1216 164 1224
rect 396 1516 404 1524
rect 540 1536 548 1544
rect 588 1836 596 1844
rect 620 1836 628 1844
rect 636 1836 644 1844
rect 732 1936 740 1944
rect 780 1936 788 1944
rect 844 2016 852 2024
rect 828 1916 836 1924
rect 668 1836 676 1844
rect 652 1816 660 1824
rect 684 1816 692 1824
rect 700 1816 708 1824
rect 620 1796 628 1804
rect 636 1796 644 1804
rect 604 1776 612 1784
rect 748 1896 756 1904
rect 796 1876 804 1884
rect 844 1876 852 1884
rect 764 1856 772 1864
rect 716 1796 724 1804
rect 668 1756 676 1764
rect 716 1756 724 1764
rect 1068 2276 1076 2284
rect 1036 2216 1044 2224
rect 1084 2196 1092 2204
rect 1020 2156 1028 2164
rect 924 2136 932 2144
rect 1020 2136 1028 2144
rect 892 2096 900 2104
rect 876 2036 884 2044
rect 892 2016 900 2024
rect 972 2116 980 2124
rect 940 2016 948 2024
rect 1084 2116 1092 2124
rect 1148 2476 1156 2484
rect 1132 2456 1140 2464
rect 1116 2296 1124 2304
rect 1212 2556 1220 2564
rect 1276 2636 1284 2644
rect 1388 2776 1396 2784
rect 1564 3856 1572 3864
rect 1516 3756 1524 3764
rect 1564 3736 1572 3744
rect 1516 3716 1524 3724
rect 1532 3616 1540 3624
rect 1740 4096 1748 4104
rect 1692 4056 1700 4064
rect 1692 4036 1700 4044
rect 1820 4336 1828 4344
rect 1804 4236 1812 4244
rect 1948 4616 1956 4624
rect 1996 4616 2004 4624
rect 2076 4576 2084 4584
rect 1916 4516 1924 4524
rect 2044 4496 2052 4504
rect 1996 4436 2004 4444
rect 1900 4356 1908 4364
rect 1932 4356 1940 4364
rect 1916 4296 1924 4304
rect 1980 4296 1988 4304
rect 1996 4276 2004 4284
rect 1900 4256 1908 4264
rect 1980 4256 1988 4264
rect 1884 4176 1892 4184
rect 1788 4116 1796 4124
rect 1772 4076 1780 4084
rect 1756 4056 1764 4064
rect 1804 4056 1812 4064
rect 1820 4056 1828 4064
rect 1788 4036 1796 4044
rect 1660 4016 1668 4024
rect 1692 3976 1700 3984
rect 1612 3836 1620 3844
rect 1660 3756 1668 3764
rect 1756 3976 1764 3984
rect 1868 4096 1876 4104
rect 1916 4176 1924 4184
rect 1852 4056 1860 4064
rect 1884 4056 1892 4064
rect 1900 4056 1908 4064
rect 1820 4036 1828 4044
rect 1836 4036 1844 4044
rect 1900 3976 1908 3984
rect 1772 3856 1780 3864
rect 1820 3876 1828 3884
rect 1708 3836 1716 3844
rect 1740 3836 1748 3844
rect 1708 3776 1716 3784
rect 1740 3776 1748 3784
rect 1612 3736 1620 3744
rect 1660 3716 1668 3724
rect 1676 3716 1684 3724
rect 1612 3696 1620 3704
rect 1596 3676 1604 3684
rect 1580 3656 1588 3664
rect 1612 3656 1620 3664
rect 1577 3606 1585 3614
rect 1587 3606 1595 3614
rect 1597 3606 1605 3614
rect 1607 3606 1615 3614
rect 1612 3576 1620 3584
rect 1548 3536 1556 3544
rect 1596 3536 1604 3544
rect 1532 3516 1540 3524
rect 1532 3496 1540 3504
rect 1580 3496 1588 3504
rect 1516 3456 1524 3464
rect 1532 3456 1540 3464
rect 1500 3396 1508 3404
rect 1452 3296 1460 3304
rect 1420 3256 1428 3264
rect 1436 3256 1444 3264
rect 1436 3016 1444 3024
rect 1436 2876 1444 2884
rect 1420 2856 1428 2864
rect 1308 2556 1316 2564
rect 1388 2676 1396 2684
rect 1420 2676 1428 2684
rect 1468 3196 1476 3204
rect 1532 3356 1540 3364
rect 1532 3336 1540 3344
rect 1500 3316 1508 3324
rect 1516 3316 1524 3324
rect 1484 3176 1492 3184
rect 1516 3196 1524 3204
rect 1564 3396 1572 3404
rect 1564 3356 1572 3364
rect 1548 3256 1556 3264
rect 1628 3556 1636 3564
rect 1612 3476 1620 3484
rect 1660 3496 1668 3504
rect 1596 3356 1604 3364
rect 1644 3396 1652 3404
rect 1580 3316 1588 3324
rect 1577 3206 1585 3214
rect 1587 3206 1595 3214
rect 1597 3206 1605 3214
rect 1607 3206 1615 3214
rect 1724 3736 1732 3744
rect 1724 3696 1732 3704
rect 1900 3876 1908 3884
rect 1884 3796 1892 3804
rect 1932 4116 1940 4124
rect 1964 4116 1972 4124
rect 1980 4116 1988 4124
rect 1948 4036 1956 4044
rect 1980 4096 1988 4104
rect 1980 4016 1988 4024
rect 1964 3876 1972 3884
rect 2028 3976 2036 3984
rect 2092 4376 2100 4384
rect 2124 4316 2132 4324
rect 2204 4516 2212 4524
rect 2172 4336 2180 4344
rect 2172 4316 2180 4324
rect 2236 4316 2244 4324
rect 2204 4276 2212 4284
rect 2460 4616 2468 4624
rect 2284 4576 2292 4584
rect 2396 4576 2404 4584
rect 2300 4536 2308 4544
rect 2444 4536 2452 4544
rect 2316 4516 2324 4524
rect 2300 4496 2308 4504
rect 2364 4496 2372 4504
rect 2268 4436 2276 4444
rect 2156 4096 2164 4104
rect 2124 4036 2132 4044
rect 2092 4016 2100 4024
rect 2076 3996 2084 4004
rect 2012 3916 2020 3924
rect 2060 3916 2068 3924
rect 1996 3876 2004 3884
rect 2108 3876 2116 3884
rect 1980 3836 1988 3844
rect 1916 3796 1924 3804
rect 1980 3796 1988 3804
rect 1852 3736 1860 3744
rect 1884 3736 1892 3744
rect 1708 3676 1716 3684
rect 1740 3676 1748 3684
rect 1692 3576 1700 3584
rect 1692 3556 1700 3564
rect 1692 3536 1700 3544
rect 1692 3496 1700 3504
rect 1772 3536 1780 3544
rect 1724 3456 1732 3464
rect 1804 3456 1812 3464
rect 1788 3436 1796 3444
rect 1708 3396 1716 3404
rect 1708 3356 1716 3364
rect 1852 3696 1860 3704
rect 1868 3696 1876 3704
rect 1836 3576 1844 3584
rect 1852 3576 1860 3584
rect 1884 3676 1892 3684
rect 1916 3756 1924 3764
rect 2060 3856 2068 3864
rect 2092 3856 2100 3864
rect 2108 3836 2116 3844
rect 2028 3816 2036 3824
rect 2220 4076 2228 4084
rect 2204 3956 2212 3964
rect 2252 4196 2260 4204
rect 2140 3916 2148 3924
rect 2140 3876 2148 3884
rect 2076 3776 2084 3784
rect 1932 3736 1940 3744
rect 2012 3736 2020 3744
rect 1916 3696 1924 3704
rect 1900 3616 1908 3624
rect 1884 3536 1892 3544
rect 1916 3536 1924 3544
rect 1836 3436 1844 3444
rect 1820 3396 1828 3404
rect 1836 3396 1844 3404
rect 1820 3376 1828 3384
rect 1676 3296 1684 3304
rect 1660 3256 1668 3264
rect 1692 3216 1700 3224
rect 1660 3196 1668 3204
rect 1532 3136 1540 3144
rect 1580 3136 1588 3144
rect 1500 3116 1508 3124
rect 1548 3116 1556 3124
rect 1564 3116 1572 3124
rect 1516 3096 1524 3104
rect 1564 3096 1572 3104
rect 1548 3076 1556 3084
rect 1468 3056 1476 3064
rect 1500 3056 1508 3064
rect 1532 3056 1540 3064
rect 1484 2896 1492 2904
rect 1500 2896 1508 2904
rect 1452 2796 1460 2804
rect 1452 2776 1460 2784
rect 1372 2656 1380 2664
rect 1372 2636 1380 2644
rect 1404 2636 1412 2644
rect 1324 2536 1332 2544
rect 1356 2536 1364 2544
rect 1388 2576 1396 2584
rect 1404 2536 1412 2544
rect 1260 2516 1268 2524
rect 1276 2516 1284 2524
rect 1388 2516 1396 2524
rect 1196 2496 1204 2504
rect 1244 2496 1252 2504
rect 1388 2476 1396 2484
rect 1404 2476 1412 2484
rect 1308 2456 1316 2464
rect 1340 2456 1348 2464
rect 1372 2456 1380 2464
rect 1420 2456 1428 2464
rect 1404 2396 1412 2404
rect 1420 2396 1428 2404
rect 1196 2336 1204 2344
rect 1164 2276 1172 2284
rect 1116 2136 1124 2144
rect 1148 2136 1156 2144
rect 1212 2296 1220 2304
rect 1212 2196 1220 2204
rect 1180 2136 1188 2144
rect 1324 2316 1332 2324
rect 1388 2316 1396 2324
rect 1404 2316 1412 2324
rect 1276 2276 1284 2284
rect 1324 2276 1332 2284
rect 1356 2276 1364 2284
rect 1260 2196 1268 2204
rect 1260 2176 1268 2184
rect 1324 2176 1332 2184
rect 1420 2276 1428 2284
rect 1404 2176 1412 2184
rect 1468 2676 1476 2684
rect 1484 2676 1492 2684
rect 1596 3096 1604 3104
rect 1580 3016 1588 3024
rect 1644 3116 1652 3124
rect 1756 3316 1764 3324
rect 1724 3256 1732 3264
rect 1724 3216 1732 3224
rect 1692 3176 1700 3184
rect 1708 3176 1716 3184
rect 1708 3116 1716 3124
rect 1660 3076 1668 3084
rect 1612 3056 1620 3064
rect 1612 2956 1620 2964
rect 1532 2916 1540 2924
rect 1532 2896 1540 2904
rect 1516 2796 1524 2804
rect 1596 2916 1604 2924
rect 1564 2896 1572 2904
rect 1644 3056 1652 3064
rect 1692 3056 1700 3064
rect 1820 3256 1828 3264
rect 1788 3216 1796 3224
rect 1868 3396 1876 3404
rect 1852 3356 1860 3364
rect 2028 3716 2036 3724
rect 2060 3716 2068 3724
rect 1964 3696 1972 3704
rect 1948 3556 1956 3564
rect 1932 3516 1940 3524
rect 2012 3616 2020 3624
rect 1996 3536 2004 3544
rect 1900 3436 1908 3444
rect 1900 3396 1908 3404
rect 1948 3476 1956 3484
rect 1932 3356 1940 3364
rect 1980 3356 1988 3364
rect 1884 3316 1892 3324
rect 1900 3256 1908 3264
rect 1932 3256 1940 3264
rect 1964 3256 1972 3264
rect 1916 3236 1924 3244
rect 1900 3176 1908 3184
rect 1788 3136 1796 3144
rect 1820 3136 1828 3144
rect 1868 3136 1876 3144
rect 1900 3136 1908 3144
rect 1868 3116 1876 3124
rect 1884 3116 1892 3124
rect 1740 3096 1748 3104
rect 1756 3076 1764 3084
rect 1740 3056 1748 3064
rect 1660 3036 1668 3044
rect 1708 3036 1716 3044
rect 1756 3016 1764 3024
rect 1676 2956 1684 2964
rect 1724 2956 1732 2964
rect 1612 2856 1620 2864
rect 1628 2856 1636 2864
rect 1548 2816 1556 2824
rect 1577 2806 1585 2814
rect 1587 2806 1595 2814
rect 1597 2806 1605 2814
rect 1607 2806 1615 2814
rect 1532 2756 1540 2764
rect 1516 2736 1524 2744
rect 1484 2656 1492 2664
rect 1500 2656 1508 2664
rect 1468 2636 1476 2644
rect 1500 2636 1508 2644
rect 1452 2476 1460 2484
rect 1452 2456 1460 2464
rect 1452 2416 1460 2424
rect 1436 2256 1444 2264
rect 1452 2236 1460 2244
rect 1372 2136 1380 2144
rect 1388 2136 1396 2144
rect 1020 2076 1028 2084
rect 988 2056 996 2064
rect 972 1996 980 2004
rect 908 1976 916 1984
rect 972 1956 980 1964
rect 892 1896 900 1904
rect 860 1776 868 1784
rect 828 1756 836 1764
rect 764 1736 772 1744
rect 588 1716 596 1724
rect 684 1716 692 1724
rect 748 1716 756 1724
rect 732 1676 740 1684
rect 716 1656 724 1664
rect 668 1576 676 1584
rect 572 1516 580 1524
rect 428 1496 436 1504
rect 524 1496 532 1504
rect 412 1456 420 1464
rect 364 1276 372 1284
rect 300 1236 308 1244
rect 124 1176 132 1184
rect 284 1176 292 1184
rect 284 1156 292 1164
rect 12 1116 20 1124
rect 220 1116 228 1124
rect 204 1096 212 1104
rect 76 1076 84 1084
rect 476 1356 484 1364
rect 412 1336 420 1344
rect 444 1316 452 1324
rect 412 1156 420 1164
rect 380 1076 388 1084
rect 44 1056 52 1064
rect 76 1056 84 1064
rect 268 1056 276 1064
rect 76 1016 84 1024
rect 92 1016 100 1024
rect 172 1036 180 1044
rect 316 1036 324 1044
rect 348 1036 356 1044
rect 332 996 340 1004
rect 124 976 132 984
rect 204 976 212 984
rect 140 956 148 964
rect 268 956 276 964
rect 364 956 372 964
rect 12 936 20 944
rect 188 936 196 944
rect 252 936 260 944
rect 300 936 308 944
rect 204 916 212 924
rect 60 736 68 744
rect 188 876 196 884
rect 252 856 260 864
rect 44 676 52 684
rect 124 676 132 684
rect 220 676 228 684
rect 12 656 20 664
rect 316 916 324 924
rect 316 816 324 824
rect 348 816 356 824
rect 332 796 340 804
rect 396 936 404 944
rect 572 1436 580 1444
rect 700 1496 708 1504
rect 604 1436 612 1444
rect 604 1396 612 1404
rect 652 1356 660 1364
rect 780 1676 788 1684
rect 748 1576 756 1584
rect 764 1576 772 1584
rect 812 1716 820 1724
rect 860 1716 868 1724
rect 796 1656 804 1664
rect 828 1656 836 1664
rect 780 1556 788 1564
rect 812 1556 820 1564
rect 732 1516 740 1524
rect 748 1516 756 1524
rect 748 1496 756 1504
rect 796 1476 804 1484
rect 700 1436 708 1444
rect 780 1436 788 1444
rect 764 1416 772 1424
rect 780 1416 788 1424
rect 748 1356 756 1364
rect 764 1356 772 1364
rect 508 1336 516 1344
rect 524 1336 532 1344
rect 588 1336 596 1344
rect 620 1336 628 1344
rect 556 1216 564 1224
rect 572 1176 580 1184
rect 492 1136 500 1144
rect 588 1136 596 1144
rect 460 1096 468 1104
rect 428 1076 436 1084
rect 460 1076 468 1084
rect 444 976 452 984
rect 428 816 436 824
rect 364 796 372 804
rect 444 716 452 724
rect 444 696 452 704
rect 348 676 356 684
rect 60 656 68 664
rect 204 656 212 664
rect 108 616 116 624
rect 172 556 180 564
rect 252 516 260 524
rect 140 496 148 504
rect 76 296 84 304
rect 108 296 116 304
rect 220 276 228 284
rect 188 256 196 264
rect 348 636 356 644
rect 380 596 388 604
rect 428 636 436 644
rect 492 1056 500 1064
rect 476 936 484 944
rect 476 916 484 924
rect 476 896 484 904
rect 524 1096 532 1104
rect 572 1096 580 1104
rect 588 1096 596 1104
rect 604 1096 612 1104
rect 572 1076 580 1084
rect 556 1056 564 1064
rect 620 1056 628 1064
rect 636 1056 644 1064
rect 572 1016 580 1024
rect 604 1016 612 1024
rect 620 996 628 1004
rect 556 956 564 964
rect 524 936 532 944
rect 508 856 516 864
rect 492 816 500 824
rect 508 816 516 824
rect 700 1256 708 1264
rect 668 1156 676 1164
rect 684 1156 692 1164
rect 764 1296 772 1304
rect 716 1236 724 1244
rect 732 1196 740 1204
rect 716 1176 724 1184
rect 700 1136 708 1144
rect 668 1056 676 1064
rect 652 916 660 924
rect 732 1156 740 1164
rect 748 1136 756 1144
rect 764 1136 772 1144
rect 732 1116 740 1124
rect 716 1056 724 1064
rect 844 1516 852 1524
rect 828 1476 836 1484
rect 844 1456 852 1464
rect 972 1876 980 1884
rect 940 1756 948 1764
rect 892 1656 900 1664
rect 1020 1936 1028 1944
rect 1004 1876 1012 1884
rect 1132 2116 1140 2124
rect 1164 2116 1172 2124
rect 1228 2116 1236 2124
rect 1324 2116 1332 2124
rect 1100 2076 1108 2084
rect 1148 2076 1156 2084
rect 1164 2076 1172 2084
rect 1196 2076 1204 2084
rect 1212 2076 1220 2084
rect 1068 1996 1076 2004
rect 1084 1996 1092 2004
rect 1148 1996 1156 2004
rect 1068 1956 1076 1964
rect 1084 1956 1092 1964
rect 1068 1876 1076 1884
rect 1036 1776 1044 1784
rect 1212 2016 1220 2024
rect 1132 1916 1140 1924
rect 1100 1896 1108 1904
rect 1164 1936 1172 1944
rect 1180 1916 1188 1924
rect 1100 1876 1108 1884
rect 1148 1876 1156 1884
rect 1100 1856 1108 1864
rect 1084 1816 1092 1824
rect 1132 1816 1140 1824
rect 1068 1776 1076 1784
rect 1100 1776 1108 1784
rect 1052 1736 1060 1744
rect 1020 1716 1028 1724
rect 1036 1696 1044 1704
rect 1036 1656 1044 1664
rect 876 1616 884 1624
rect 956 1616 964 1624
rect 1052 1636 1060 1644
rect 1244 1996 1252 2004
rect 1276 1996 1284 2004
rect 1244 1956 1252 1964
rect 1276 1956 1284 1964
rect 1372 2076 1380 2084
rect 1452 2156 1460 2164
rect 1516 2576 1524 2584
rect 1660 2856 1668 2864
rect 1676 2856 1684 2864
rect 1548 2736 1556 2744
rect 1564 2736 1572 2744
rect 1644 2736 1652 2744
rect 1564 2696 1572 2704
rect 1548 2676 1556 2684
rect 1596 2656 1604 2664
rect 1596 2636 1604 2644
rect 1612 2636 1620 2644
rect 1564 2576 1572 2584
rect 1564 2556 1572 2564
rect 1596 2556 1604 2564
rect 1500 2476 1508 2484
rect 1532 2476 1540 2484
rect 1516 2436 1524 2444
rect 1484 2396 1492 2404
rect 1516 2376 1524 2384
rect 1532 2376 1540 2384
rect 1500 2356 1508 2364
rect 1484 2316 1492 2324
rect 1516 2316 1524 2324
rect 1676 2816 1684 2824
rect 1788 3056 1796 3064
rect 1884 3076 1892 3084
rect 1852 3056 1860 3064
rect 1820 3036 1828 3044
rect 1836 3036 1844 3044
rect 1756 2896 1764 2904
rect 1772 2876 1780 2884
rect 1708 2856 1716 2864
rect 1692 2796 1700 2804
rect 1676 2756 1684 2764
rect 1676 2716 1684 2724
rect 1692 2676 1700 2684
rect 1692 2656 1700 2664
rect 1756 2776 1764 2784
rect 1868 2996 1876 3004
rect 1820 2916 1828 2924
rect 1868 2916 1876 2924
rect 1932 3216 1940 3224
rect 1932 3136 1940 3144
rect 1964 3136 1972 3144
rect 2060 3616 2068 3624
rect 2028 3536 2036 3544
rect 2012 3516 2020 3524
rect 2044 3516 2052 3524
rect 2028 3476 2036 3484
rect 2108 3716 2116 3724
rect 2108 3696 2116 3704
rect 2108 3656 2116 3664
rect 2108 3596 2116 3604
rect 2092 3556 2100 3564
rect 2076 3516 2084 3524
rect 2076 3496 2084 3504
rect 2156 3856 2164 3864
rect 2188 3856 2196 3864
rect 2220 3816 2228 3824
rect 2188 3776 2196 3784
rect 2156 3716 2164 3724
rect 2172 3656 2180 3664
rect 2156 3556 2164 3564
rect 2108 3476 2116 3484
rect 2060 3436 2068 3444
rect 2204 3576 2212 3584
rect 2172 3476 2180 3484
rect 2044 3356 2052 3364
rect 2124 3416 2132 3424
rect 2076 3396 2084 3404
rect 2092 3356 2100 3364
rect 2108 3356 2116 3364
rect 2156 3356 2164 3364
rect 2204 3496 2212 3504
rect 2204 3456 2212 3464
rect 2044 3296 2052 3304
rect 2108 3276 2116 3284
rect 2060 3256 2068 3264
rect 2012 3196 2020 3204
rect 1996 3136 2004 3144
rect 2028 3136 2036 3144
rect 1980 3116 1988 3124
rect 1964 3096 1972 3104
rect 2092 3236 2100 3244
rect 2060 3116 2068 3124
rect 2060 3096 2068 3104
rect 1932 3076 1940 3084
rect 1900 2996 1908 3004
rect 1964 3056 1972 3064
rect 1932 2956 1940 2964
rect 2044 3056 2052 3064
rect 2028 3036 2036 3044
rect 2044 3036 2052 3044
rect 1980 3016 1988 3024
rect 1996 3016 2004 3024
rect 2044 2996 2052 3004
rect 1900 2916 1908 2924
rect 1852 2876 1860 2884
rect 1884 2876 1892 2884
rect 1836 2856 1844 2864
rect 1788 2816 1796 2824
rect 1804 2816 1812 2824
rect 1804 2796 1812 2804
rect 1788 2756 1796 2764
rect 1804 2756 1812 2764
rect 1772 2736 1780 2744
rect 1756 2716 1764 2724
rect 1820 2736 1828 2744
rect 1820 2716 1828 2724
rect 1708 2636 1716 2644
rect 1724 2636 1732 2644
rect 1660 2556 1668 2564
rect 1692 2556 1700 2564
rect 1628 2476 1636 2484
rect 1772 2676 1780 2684
rect 1804 2656 1812 2664
rect 1804 2636 1812 2644
rect 1820 2636 1828 2644
rect 1676 2536 1684 2544
rect 1756 2536 1764 2544
rect 1660 2416 1668 2424
rect 1577 2406 1585 2414
rect 1587 2406 1595 2414
rect 1597 2406 1605 2414
rect 1607 2406 1615 2414
rect 1644 2396 1652 2404
rect 1580 2356 1588 2364
rect 1548 2276 1556 2284
rect 1500 2156 1508 2164
rect 1772 2516 1780 2524
rect 1724 2436 1732 2444
rect 1756 2436 1764 2444
rect 1708 2416 1716 2424
rect 1724 2356 1732 2364
rect 1708 2316 1716 2324
rect 1692 2276 1700 2284
rect 1660 2256 1668 2264
rect 1676 2256 1684 2264
rect 1724 2256 1732 2264
rect 1756 2276 1764 2284
rect 1724 2156 1732 2164
rect 1564 2136 1572 2144
rect 1644 2136 1652 2144
rect 1708 2136 1716 2144
rect 1724 2136 1732 2144
rect 1676 2116 1684 2124
rect 1532 2076 1540 2084
rect 1596 2096 1604 2104
rect 1660 2096 1668 2104
rect 1340 2016 1348 2024
rect 1404 2016 1412 2024
rect 1468 2016 1476 2024
rect 1577 2006 1585 2014
rect 1587 2006 1595 2014
rect 1597 2006 1605 2014
rect 1607 2006 1615 2014
rect 1340 1996 1348 2004
rect 1356 1996 1364 2004
rect 1372 1996 1380 2004
rect 1484 1996 1492 2004
rect 1516 1996 1524 2004
rect 1324 1956 1332 1964
rect 1244 1916 1252 1924
rect 1692 2056 1700 2064
rect 1660 2016 1668 2024
rect 1660 1996 1668 2004
rect 1676 1956 1684 1964
rect 1644 1936 1652 1944
rect 1612 1916 1620 1924
rect 1260 1836 1268 1844
rect 1228 1816 1236 1824
rect 1244 1816 1252 1824
rect 1308 1876 1316 1884
rect 1324 1876 1332 1884
rect 1292 1856 1300 1864
rect 1196 1796 1204 1804
rect 1212 1796 1220 1804
rect 1164 1736 1172 1744
rect 1068 1616 1076 1624
rect 1148 1616 1156 1624
rect 1036 1556 1044 1564
rect 988 1536 996 1544
rect 940 1516 948 1524
rect 1052 1516 1060 1524
rect 1084 1516 1092 1524
rect 1132 1536 1140 1544
rect 876 1496 884 1504
rect 988 1496 996 1504
rect 1020 1496 1028 1504
rect 1052 1496 1060 1504
rect 1100 1496 1108 1504
rect 876 1476 884 1484
rect 892 1476 900 1484
rect 860 1436 868 1444
rect 828 1416 836 1424
rect 860 1416 868 1424
rect 876 1416 884 1424
rect 796 1316 804 1324
rect 780 1116 788 1124
rect 732 976 740 984
rect 700 936 708 944
rect 748 936 756 944
rect 700 916 708 924
rect 556 876 564 884
rect 668 876 676 884
rect 684 876 692 884
rect 524 716 532 724
rect 540 716 548 724
rect 492 696 500 704
rect 636 856 644 864
rect 668 856 676 864
rect 748 836 756 844
rect 748 816 756 824
rect 812 1216 820 1224
rect 812 1136 820 1144
rect 844 1136 852 1144
rect 844 1056 852 1064
rect 988 1456 996 1464
rect 940 1376 948 1384
rect 956 1376 964 1384
rect 972 1376 980 1384
rect 1020 1416 1028 1424
rect 1036 1416 1044 1424
rect 1132 1476 1140 1484
rect 1148 1476 1156 1484
rect 1052 1396 1060 1404
rect 1116 1416 1124 1424
rect 1020 1336 1028 1344
rect 1036 1336 1044 1344
rect 1084 1336 1092 1344
rect 1100 1336 1108 1344
rect 876 1316 884 1324
rect 892 1316 900 1324
rect 956 1316 964 1324
rect 892 1296 900 1304
rect 924 1296 932 1304
rect 1068 1296 1076 1304
rect 1084 1296 1092 1304
rect 1052 1256 1060 1264
rect 924 1196 932 1204
rect 972 1196 980 1204
rect 924 1176 932 1184
rect 956 1116 964 1124
rect 1004 1216 1012 1224
rect 1036 1216 1044 1224
rect 876 1056 884 1064
rect 828 996 836 1004
rect 796 896 804 904
rect 828 896 836 904
rect 780 816 788 824
rect 716 776 724 784
rect 716 736 724 744
rect 620 716 628 724
rect 636 716 644 724
rect 684 716 692 724
rect 764 796 772 804
rect 764 776 772 784
rect 780 716 788 724
rect 812 816 820 824
rect 860 996 868 1004
rect 860 956 868 964
rect 892 996 900 1004
rect 876 936 884 944
rect 940 1036 948 1044
rect 988 1016 996 1024
rect 924 996 932 1004
rect 956 996 964 1004
rect 972 996 980 1004
rect 1132 1396 1140 1404
rect 1276 1796 1284 1804
rect 1244 1736 1252 1744
rect 1244 1616 1252 1624
rect 1244 1596 1252 1604
rect 1228 1536 1236 1544
rect 1340 1816 1348 1824
rect 1356 1816 1364 1824
rect 1292 1776 1300 1784
rect 1388 1816 1396 1824
rect 1372 1796 1380 1804
rect 1740 2116 1748 2124
rect 1756 2096 1764 2104
rect 1788 2356 1796 2364
rect 1788 2316 1796 2324
rect 1788 2256 1796 2264
rect 1932 2876 1940 2884
rect 1916 2716 1924 2724
rect 1948 2816 1956 2824
rect 1852 2696 1860 2704
rect 1884 2696 1892 2704
rect 1852 2676 1860 2684
rect 1820 2616 1828 2624
rect 1836 2616 1844 2624
rect 1916 2676 1924 2684
rect 1948 2676 1956 2684
rect 1964 2676 1972 2684
rect 1900 2656 1908 2664
rect 1884 2636 1892 2644
rect 1820 2536 1828 2544
rect 1948 2616 1956 2624
rect 1852 2556 1860 2564
rect 1868 2556 1876 2564
rect 1900 2556 1908 2564
rect 1916 2556 1924 2564
rect 1884 2536 1892 2544
rect 1932 2536 1940 2544
rect 1852 2476 1860 2484
rect 1852 2436 1860 2444
rect 1820 2376 1828 2384
rect 1884 2436 1892 2444
rect 1964 2576 1972 2584
rect 1948 2496 1956 2504
rect 1932 2416 1940 2424
rect 1884 2376 1892 2384
rect 1948 2376 1956 2384
rect 1852 2356 1860 2364
rect 1868 2356 1876 2364
rect 1884 2316 1892 2324
rect 1900 2316 1908 2324
rect 1932 2316 1940 2324
rect 1820 2276 1828 2284
rect 2028 2956 2036 2964
rect 1996 2876 2004 2884
rect 1996 2836 2004 2844
rect 2012 2836 2020 2844
rect 1996 2796 2004 2804
rect 1996 2676 2004 2684
rect 2044 2836 2052 2844
rect 2076 3056 2084 3064
rect 2092 3056 2100 3064
rect 2076 2996 2084 3004
rect 2156 3296 2164 3304
rect 2140 3256 2148 3264
rect 2140 3216 2148 3224
rect 2156 3156 2164 3164
rect 2124 3116 2132 3124
rect 2204 3336 2212 3344
rect 2188 3316 2196 3324
rect 2204 3316 2212 3324
rect 2252 3916 2260 3924
rect 2252 3716 2260 3724
rect 2332 4436 2340 4444
rect 2396 4436 2404 4444
rect 2300 4416 2308 4424
rect 2284 4376 2292 4384
rect 2332 4376 2340 4384
rect 2284 4316 2292 4324
rect 2300 4316 2308 4324
rect 2380 4316 2388 4324
rect 2300 4296 2308 4304
rect 2460 4376 2468 4384
rect 2428 4316 2436 4324
rect 2316 4276 2324 4284
rect 2380 4196 2388 4204
rect 2284 4176 2292 4184
rect 2284 4116 2292 4124
rect 2412 4216 2420 4224
rect 2396 4096 2404 4104
rect 2300 4036 2308 4044
rect 2380 3936 2388 3944
rect 2492 4176 2500 4184
rect 2748 4616 2756 4624
rect 2908 4616 2916 4624
rect 3084 4616 3092 4624
rect 3244 4616 3252 4624
rect 3308 4616 3316 4624
rect 3500 4616 3508 4624
rect 3516 4616 3524 4624
rect 2860 4576 2868 4584
rect 2572 4556 2580 4564
rect 2732 4556 2740 4564
rect 2924 4556 2932 4564
rect 3052 4556 3060 4564
rect 3068 4556 3076 4564
rect 2684 4536 2692 4544
rect 2780 4536 2788 4544
rect 2668 4516 2676 4524
rect 2716 4516 2724 4524
rect 2780 4516 2788 4524
rect 2812 4516 2820 4524
rect 2892 4518 2900 4524
rect 2892 4516 2900 4518
rect 2892 4496 2900 4504
rect 2652 4376 2660 4384
rect 2732 4376 2740 4384
rect 2684 4356 2692 4364
rect 2556 4336 2564 4344
rect 2524 4296 2532 4304
rect 2540 4296 2548 4304
rect 2908 4336 2916 4344
rect 2956 4536 2964 4544
rect 3020 4496 3028 4504
rect 2828 4316 2836 4324
rect 2924 4316 2932 4324
rect 2956 4316 2964 4324
rect 2700 4296 2708 4304
rect 2748 4296 2756 4304
rect 2844 4296 2852 4304
rect 2876 4296 2884 4304
rect 2940 4296 2948 4304
rect 2700 4256 2708 4264
rect 2524 4236 2532 4244
rect 2556 4116 2564 4124
rect 2492 4096 2500 4104
rect 2524 4096 2532 4104
rect 2540 4096 2548 4104
rect 2604 4096 2612 4104
rect 2620 4096 2628 4104
rect 2444 4016 2452 4024
rect 2428 3936 2436 3944
rect 2332 3916 2340 3924
rect 2316 3896 2324 3904
rect 2284 3836 2292 3844
rect 2236 3596 2244 3604
rect 2236 3476 2244 3484
rect 2396 3896 2404 3904
rect 2428 3896 2436 3904
rect 2396 3876 2404 3884
rect 2428 3876 2436 3884
rect 2412 3856 2420 3864
rect 2348 3836 2356 3844
rect 2396 3836 2404 3844
rect 2364 3796 2372 3804
rect 2460 3976 2468 3984
rect 2588 4076 2596 4084
rect 2668 4076 2676 4084
rect 2556 4036 2564 4044
rect 2540 3996 2548 4004
rect 2556 3996 2564 4004
rect 2444 3856 2452 3864
rect 2492 3956 2500 3964
rect 2492 3916 2500 3924
rect 2476 3876 2484 3884
rect 2524 3856 2532 3864
rect 2572 3876 2580 3884
rect 2588 3876 2596 3884
rect 2556 3856 2564 3864
rect 2348 3736 2356 3744
rect 2364 3736 2372 3744
rect 2460 3736 2468 3744
rect 2540 3736 2548 3744
rect 2332 3656 2340 3664
rect 2300 3616 2308 3624
rect 2204 3216 2212 3224
rect 2204 3096 2212 3104
rect 2284 3456 2292 3464
rect 2332 3536 2340 3544
rect 2316 3456 2324 3464
rect 2332 3456 2340 3464
rect 2268 3416 2276 3424
rect 2300 3416 2308 3424
rect 2300 3396 2308 3404
rect 2444 3716 2452 3724
rect 2412 3696 2420 3704
rect 2428 3676 2436 3684
rect 2380 3576 2388 3584
rect 2460 3696 2468 3704
rect 2508 3696 2516 3704
rect 2492 3676 2500 3684
rect 2476 3616 2484 3624
rect 2460 3596 2468 3604
rect 2396 3536 2404 3544
rect 2428 3536 2436 3544
rect 2444 3536 2452 3544
rect 2380 3516 2388 3524
rect 2428 3496 2436 3504
rect 2460 3496 2468 3504
rect 2428 3476 2436 3484
rect 2444 3476 2452 3484
rect 2348 3396 2356 3404
rect 2380 3396 2388 3404
rect 2348 3376 2356 3384
rect 2364 3376 2372 3384
rect 2364 3356 2372 3364
rect 2252 3316 2260 3324
rect 2268 3316 2276 3324
rect 2316 3316 2324 3324
rect 2348 3316 2356 3324
rect 2284 3256 2292 3264
rect 2332 3256 2340 3264
rect 2364 3256 2372 3264
rect 2412 3316 2420 3324
rect 2428 3316 2436 3324
rect 2380 3176 2388 3184
rect 2396 3176 2404 3184
rect 2284 3156 2292 3164
rect 2316 3156 2324 3164
rect 2268 3116 2276 3124
rect 2172 3056 2180 3064
rect 2140 2996 2148 3004
rect 2268 3076 2276 3084
rect 2252 3056 2260 3064
rect 2284 3056 2292 3064
rect 2252 3036 2260 3044
rect 2236 3016 2244 3024
rect 2092 2896 2100 2904
rect 2108 2876 2116 2884
rect 2108 2836 2116 2844
rect 2188 2996 2196 3004
rect 2204 2996 2212 3004
rect 2268 3016 2276 3024
rect 2188 2956 2196 2964
rect 2204 2956 2212 2964
rect 2252 2956 2260 2964
rect 2156 2896 2164 2904
rect 2172 2896 2180 2904
rect 2188 2876 2196 2884
rect 2140 2856 2148 2864
rect 2156 2856 2164 2864
rect 2124 2816 2132 2824
rect 2268 2936 2276 2944
rect 2220 2876 2228 2884
rect 2156 2816 2164 2824
rect 2204 2816 2212 2824
rect 2188 2776 2196 2784
rect 2076 2696 2084 2704
rect 2044 2656 2052 2664
rect 2028 2616 2036 2624
rect 2012 2576 2020 2584
rect 2044 2576 2052 2584
rect 2060 2576 2068 2584
rect 1996 2556 2004 2564
rect 2012 2556 2020 2564
rect 2092 2656 2100 2664
rect 2124 2616 2132 2624
rect 2140 2616 2148 2624
rect 1980 2536 1988 2544
rect 2012 2536 2020 2544
rect 2092 2556 2100 2564
rect 2060 2536 2068 2544
rect 1964 2336 1972 2344
rect 1836 2236 1844 2244
rect 1852 2236 1860 2244
rect 1804 2176 1812 2184
rect 1916 2216 1924 2224
rect 1884 2196 1892 2204
rect 1980 2276 1988 2284
rect 1964 2256 1972 2264
rect 1788 2096 1796 2104
rect 1756 1996 1764 2004
rect 1708 1916 1716 1924
rect 1724 1916 1732 1924
rect 1756 1916 1764 1924
rect 1468 1876 1476 1884
rect 1484 1876 1492 1884
rect 1644 1876 1652 1884
rect 1676 1896 1684 1904
rect 1724 1896 1732 1904
rect 1772 1876 1780 1884
rect 1548 1856 1556 1864
rect 1436 1816 1444 1824
rect 1420 1796 1428 1804
rect 1468 1816 1476 1824
rect 1644 1836 1652 1844
rect 1452 1796 1460 1804
rect 1484 1796 1492 1804
rect 1500 1796 1508 1804
rect 1372 1716 1380 1724
rect 1324 1696 1332 1704
rect 1340 1696 1348 1704
rect 1372 1696 1380 1704
rect 1276 1616 1284 1624
rect 1484 1716 1492 1724
rect 1468 1676 1476 1684
rect 1324 1596 1332 1604
rect 1292 1536 1300 1544
rect 1196 1516 1204 1524
rect 1260 1516 1268 1524
rect 1244 1496 1252 1504
rect 1260 1496 1268 1504
rect 1164 1336 1172 1344
rect 1116 1296 1124 1304
rect 1148 1296 1156 1304
rect 1100 1236 1108 1244
rect 1132 1236 1140 1244
rect 1116 1216 1124 1224
rect 1052 1136 1060 1144
rect 1020 1016 1028 1024
rect 940 976 948 984
rect 812 776 820 784
rect 908 756 916 764
rect 1020 976 1028 984
rect 988 956 996 964
rect 1004 956 1012 964
rect 1020 936 1028 944
rect 972 896 980 904
rect 988 896 996 904
rect 956 876 964 884
rect 940 776 948 784
rect 828 716 836 724
rect 572 676 580 684
rect 620 676 628 684
rect 476 636 484 644
rect 524 636 532 644
rect 444 616 452 624
rect 460 616 468 624
rect 412 576 420 584
rect 508 616 516 624
rect 556 616 564 624
rect 444 556 452 564
rect 604 656 612 664
rect 588 556 596 564
rect 492 536 500 544
rect 556 536 564 544
rect 572 536 580 544
rect 588 496 596 504
rect 636 556 644 564
rect 652 556 660 564
rect 620 536 628 544
rect 844 616 852 624
rect 716 576 724 584
rect 796 576 804 584
rect 652 536 660 544
rect 668 536 676 544
rect 604 476 612 484
rect 620 476 628 484
rect 636 476 644 484
rect 380 376 388 384
rect 572 356 580 364
rect 316 296 324 304
rect 460 296 468 304
rect 540 256 548 264
rect 332 196 340 204
rect 700 516 708 524
rect 732 556 740 564
rect 748 556 756 564
rect 812 556 820 564
rect 828 556 836 564
rect 748 516 756 524
rect 780 496 788 504
rect 812 496 820 504
rect 748 476 756 484
rect 764 476 772 484
rect 732 416 740 424
rect 684 296 692 304
rect 652 216 660 224
rect 764 176 772 184
rect 860 536 868 544
rect 892 676 900 684
rect 940 696 948 704
rect 956 676 964 684
rect 1084 1116 1092 1124
rect 1132 1116 1140 1124
rect 1212 1476 1220 1484
rect 1228 1476 1236 1484
rect 1228 1416 1236 1424
rect 1212 1316 1220 1324
rect 1260 1456 1268 1464
rect 1260 1336 1268 1344
rect 1212 1296 1220 1304
rect 1244 1296 1252 1304
rect 1212 1276 1220 1284
rect 1196 1256 1204 1264
rect 1180 1236 1188 1244
rect 1148 1096 1156 1104
rect 1164 1076 1172 1084
rect 1116 1056 1124 1064
rect 1116 1036 1124 1044
rect 1100 996 1108 1004
rect 1084 976 1092 984
rect 1068 956 1076 964
rect 1084 956 1092 964
rect 1052 936 1060 944
rect 1068 936 1076 944
rect 1052 816 1060 824
rect 1068 816 1076 824
rect 1036 796 1044 804
rect 1148 1056 1156 1064
rect 1132 1016 1140 1024
rect 1132 976 1140 984
rect 1116 896 1124 904
rect 1116 856 1124 864
rect 1100 796 1108 804
rect 1084 756 1092 764
rect 988 696 996 704
rect 1052 716 1060 724
rect 1020 696 1028 704
rect 1052 696 1060 704
rect 1196 1096 1204 1104
rect 1260 1196 1268 1204
rect 1292 1376 1300 1384
rect 1324 1536 1332 1544
rect 1468 1596 1476 1604
rect 1404 1516 1412 1524
rect 1420 1516 1428 1524
rect 1468 1516 1476 1524
rect 1644 1816 1652 1824
rect 1884 2116 1892 2124
rect 1948 2176 1956 2184
rect 1964 2156 1972 2164
rect 1836 2016 1844 2024
rect 1804 1996 1812 2004
rect 1804 1976 1812 1984
rect 1836 1976 1844 1984
rect 1804 1896 1812 1904
rect 1676 1836 1684 1844
rect 1772 1836 1780 1844
rect 1788 1836 1796 1844
rect 1628 1796 1636 1804
rect 1660 1796 1668 1804
rect 1692 1816 1700 1824
rect 1708 1816 1716 1824
rect 1516 1696 1524 1704
rect 1516 1676 1524 1684
rect 1532 1616 1540 1624
rect 1516 1596 1524 1604
rect 1500 1516 1508 1524
rect 1340 1436 1348 1444
rect 1324 1276 1332 1284
rect 1308 1256 1316 1264
rect 1324 1236 1332 1244
rect 1244 1136 1252 1144
rect 1260 1136 1268 1144
rect 1292 1136 1300 1144
rect 1308 1136 1316 1144
rect 1388 1456 1396 1464
rect 1420 1496 1428 1504
rect 1468 1496 1476 1504
rect 1404 1416 1412 1424
rect 1404 1356 1412 1364
rect 1372 1336 1380 1344
rect 1388 1336 1396 1344
rect 1436 1476 1444 1484
rect 1532 1516 1540 1524
rect 1644 1616 1652 1624
rect 1577 1606 1585 1614
rect 1587 1606 1595 1614
rect 1597 1606 1605 1614
rect 1607 1606 1615 1614
rect 1644 1596 1652 1604
rect 1660 1576 1668 1584
rect 1436 1356 1444 1364
rect 1452 1356 1460 1364
rect 1372 1296 1380 1304
rect 1356 1256 1364 1264
rect 1356 1236 1364 1244
rect 1244 1116 1252 1124
rect 1308 1116 1316 1124
rect 1324 1116 1332 1124
rect 1260 1036 1268 1044
rect 1292 1036 1300 1044
rect 1148 956 1156 964
rect 1244 976 1252 984
rect 1228 956 1236 964
rect 1244 936 1252 944
rect 1276 936 1284 944
rect 1132 776 1140 784
rect 1180 856 1188 864
rect 1212 876 1220 884
rect 1260 896 1268 904
rect 1196 796 1204 804
rect 1244 796 1252 804
rect 1148 756 1156 764
rect 1180 756 1188 764
rect 1116 736 1124 744
rect 1340 1016 1348 1024
rect 1436 1336 1444 1344
rect 1484 1336 1492 1344
rect 1532 1456 1540 1464
rect 1596 1496 1604 1504
rect 1596 1456 1604 1464
rect 1596 1416 1604 1424
rect 1580 1376 1588 1384
rect 1548 1336 1556 1344
rect 1564 1336 1572 1344
rect 1532 1316 1540 1324
rect 1436 1296 1444 1304
rect 1404 1276 1412 1284
rect 1436 1276 1444 1284
rect 1500 1296 1508 1304
rect 1436 1236 1444 1244
rect 1452 1236 1460 1244
rect 1468 1216 1476 1224
rect 1404 1196 1412 1204
rect 1420 1136 1428 1144
rect 1436 1136 1444 1144
rect 1388 1096 1396 1104
rect 1404 1096 1412 1104
rect 1372 1016 1380 1024
rect 1532 1276 1540 1284
rect 1644 1536 1652 1544
rect 1740 1736 1748 1744
rect 1900 2076 1908 2084
rect 1916 2076 1924 2084
rect 1868 1956 1876 1964
rect 1884 1956 1892 1964
rect 1788 1816 1796 1824
rect 1820 1816 1828 1824
rect 1836 1816 1844 1824
rect 1852 1816 1860 1824
rect 1900 1896 1908 1904
rect 1948 1976 1956 1984
rect 2220 2736 2228 2744
rect 2204 2676 2212 2684
rect 2300 3016 2308 3024
rect 2444 3296 2452 3304
rect 2492 3476 2500 3484
rect 2556 3596 2564 3604
rect 2668 3996 2676 4004
rect 2652 3976 2660 3984
rect 2636 3916 2644 3924
rect 2668 3916 2676 3924
rect 2620 3876 2628 3884
rect 2604 3856 2612 3864
rect 2652 3876 2660 3884
rect 2604 3796 2612 3804
rect 2636 3796 2644 3804
rect 2524 3576 2532 3584
rect 2636 3716 2644 3724
rect 2604 3556 2612 3564
rect 2620 3536 2628 3544
rect 2556 3516 2564 3524
rect 2540 3496 2548 3504
rect 2476 3396 2484 3404
rect 2508 3396 2516 3404
rect 2540 3376 2548 3384
rect 2524 3316 2532 3324
rect 2780 4236 2788 4244
rect 2860 4216 2868 4224
rect 2828 4156 2836 4164
rect 2812 4136 2820 4144
rect 2924 4236 2932 4244
rect 2908 4196 2916 4204
rect 2924 4196 2932 4204
rect 2860 4116 2868 4124
rect 2940 4116 2948 4124
rect 2716 4076 2724 4084
rect 2780 4076 2788 4084
rect 2812 4076 2820 4084
rect 2876 4076 2884 4084
rect 2892 4076 2900 4084
rect 2908 4076 2916 4084
rect 2764 3996 2772 4004
rect 2748 3976 2756 3984
rect 2700 3936 2708 3944
rect 2716 3936 2724 3944
rect 2684 3856 2692 3864
rect 2668 3776 2676 3784
rect 2684 3776 2692 3784
rect 2748 3876 2756 3884
rect 2716 3856 2724 3864
rect 2684 3736 2692 3744
rect 2700 3736 2708 3744
rect 2668 3716 2676 3724
rect 2668 3696 2676 3704
rect 2652 3536 2660 3544
rect 2572 3476 2580 3484
rect 2588 3476 2596 3484
rect 2604 3456 2612 3464
rect 2588 3376 2596 3384
rect 2620 3376 2628 3384
rect 2572 3336 2580 3344
rect 2492 3296 2500 3304
rect 2508 3256 2516 3264
rect 2524 3256 2532 3264
rect 2460 3216 2468 3224
rect 2492 3216 2500 3224
rect 2428 3156 2436 3164
rect 2444 3156 2452 3164
rect 2428 3136 2436 3144
rect 2364 3116 2372 3124
rect 2380 3116 2388 3124
rect 2348 3076 2356 3084
rect 2396 3076 2404 3084
rect 2364 3056 2372 3064
rect 2604 3356 2612 3364
rect 2604 3336 2612 3344
rect 2636 3336 2644 3344
rect 2604 3296 2612 3304
rect 2636 3296 2644 3304
rect 2588 3256 2596 3264
rect 2604 3256 2612 3264
rect 2604 3196 2612 3204
rect 2700 3696 2708 3704
rect 2700 3676 2708 3684
rect 2748 3756 2756 3764
rect 2732 3676 2740 3684
rect 2716 3656 2724 3664
rect 2700 3596 2708 3604
rect 2716 3596 2724 3604
rect 2684 3496 2692 3504
rect 2780 3936 2788 3944
rect 2780 3916 2788 3924
rect 2860 4056 2868 4064
rect 2876 3996 2884 4004
rect 2892 3996 2900 4004
rect 2876 3956 2884 3964
rect 2892 3896 2900 3904
rect 2972 4296 2980 4304
rect 3004 4296 3012 4304
rect 3052 4456 3060 4464
rect 2972 4256 2980 4264
rect 2988 4256 2996 4264
rect 2988 4196 2996 4204
rect 2972 4076 2980 4084
rect 3052 4256 3060 4264
rect 3036 4136 3044 4144
rect 3004 4116 3012 4124
rect 3020 4096 3028 4104
rect 2956 3936 2964 3944
rect 2780 3876 2788 3884
rect 2796 3876 2804 3884
rect 2812 3876 2820 3884
rect 2860 3876 2868 3884
rect 2908 3876 2916 3884
rect 2828 3856 2836 3864
rect 2860 3796 2868 3804
rect 2812 3756 2820 3764
rect 2828 3736 2836 3744
rect 2924 3796 2932 3804
rect 2908 3756 2916 3764
rect 3113 4606 3121 4614
rect 3123 4606 3131 4614
rect 3133 4606 3141 4614
rect 3143 4606 3151 4614
rect 3356 4556 3364 4564
rect 3260 4536 3268 4544
rect 3420 4536 3428 4544
rect 3164 4516 3172 4524
rect 3084 4496 3092 4504
rect 3100 4476 3108 4484
rect 3116 4456 3124 4464
rect 3356 4516 3364 4524
rect 3420 4516 3428 4524
rect 3372 4476 3380 4484
rect 3276 4336 3284 4344
rect 3180 4316 3188 4324
rect 3113 4206 3121 4214
rect 3123 4206 3131 4214
rect 3133 4206 3141 4214
rect 3143 4206 3151 4214
rect 3148 4156 3156 4164
rect 3084 4116 3092 4124
rect 3068 4096 3076 4104
rect 3100 4076 3108 4084
rect 3212 4276 3220 4284
rect 3228 4276 3236 4284
rect 5932 4596 5940 4604
rect 6236 4596 6244 4604
rect 4060 4576 4068 4584
rect 4092 4576 4100 4584
rect 4700 4556 4708 4564
rect 4812 4556 4820 4564
rect 4828 4556 4836 4564
rect 5356 4556 5364 4564
rect 5612 4556 5620 4564
rect 5788 4556 5796 4564
rect 3516 4536 3524 4544
rect 4204 4536 4212 4544
rect 4716 4536 4724 4544
rect 4780 4536 4788 4544
rect 4940 4536 4948 4544
rect 3532 4516 3540 4524
rect 3484 4496 3492 4504
rect 3532 4496 3540 4504
rect 3804 4496 3812 4504
rect 3452 4456 3460 4464
rect 3660 4476 3668 4484
rect 3644 4456 3652 4464
rect 3644 4416 3652 4424
rect 3548 4336 3556 4344
rect 3372 4316 3380 4324
rect 3500 4316 3508 4324
rect 3580 4316 3588 4324
rect 3612 4316 3616 4324
rect 3616 4316 3620 4324
rect 3372 4296 3380 4304
rect 3404 4296 3412 4304
rect 3292 4216 3300 4224
rect 3228 4196 3236 4204
rect 3324 4176 3332 4184
rect 3308 4156 3316 4164
rect 3276 4136 3284 4144
rect 3244 4116 3252 4124
rect 3196 4096 3204 4104
rect 3228 4096 3236 4104
rect 3116 3936 3124 3944
rect 3020 3876 3028 3884
rect 2780 3716 2788 3724
rect 2876 3716 2884 3724
rect 2908 3716 2916 3724
rect 2780 3616 2788 3624
rect 2828 3656 2836 3664
rect 2828 3616 2836 3624
rect 2796 3596 2804 3604
rect 2892 3676 2900 3684
rect 2908 3676 2916 3684
rect 2956 3676 2964 3684
rect 2972 3676 2980 3684
rect 2908 3616 2916 3624
rect 2908 3596 2916 3604
rect 2828 3556 2836 3564
rect 2876 3556 2884 3564
rect 2796 3536 2804 3544
rect 2748 3456 2756 3464
rect 2668 3436 2676 3444
rect 2732 3436 2740 3444
rect 2844 3536 2852 3544
rect 2892 3516 2900 3524
rect 2972 3656 2980 3664
rect 2972 3596 2980 3604
rect 2828 3416 2836 3424
rect 2892 3476 2900 3484
rect 2876 3456 2884 3464
rect 2972 3436 2980 3444
rect 2908 3416 2916 3424
rect 2796 3376 2804 3384
rect 2844 3376 2852 3384
rect 2668 3356 2676 3364
rect 2780 3356 2788 3364
rect 2748 3316 2756 3324
rect 2668 3296 2676 3304
rect 2716 3296 2724 3304
rect 2700 3256 2708 3264
rect 2652 3156 2660 3164
rect 2508 3136 2516 3144
rect 2540 3136 2548 3144
rect 2460 3076 2468 3084
rect 2396 3036 2404 3044
rect 2412 3036 2420 3044
rect 2444 3036 2452 3044
rect 2348 2996 2356 3004
rect 2364 2996 2372 3004
rect 2300 2956 2308 2964
rect 2316 2956 2324 2964
rect 2348 2936 2356 2944
rect 2332 2896 2340 2904
rect 2364 2896 2372 2904
rect 2380 2896 2388 2904
rect 2348 2876 2356 2884
rect 2332 2856 2340 2864
rect 2284 2836 2292 2844
rect 2284 2816 2292 2824
rect 2252 2736 2260 2744
rect 2364 2716 2372 2724
rect 2188 2656 2196 2664
rect 2172 2556 2180 2564
rect 2188 2556 2196 2564
rect 2124 2516 2132 2524
rect 2012 2476 2020 2484
rect 2028 2476 2036 2484
rect 2092 2436 2100 2444
rect 2076 2416 2084 2424
rect 2028 2356 2036 2364
rect 2108 2396 2116 2404
rect 2124 2356 2132 2364
rect 2300 2676 2308 2684
rect 2316 2676 2324 2684
rect 2236 2636 2244 2644
rect 2220 2616 2228 2624
rect 2300 2616 2308 2624
rect 2444 2916 2452 2924
rect 2460 2876 2468 2884
rect 2428 2816 2436 2824
rect 2444 2776 2452 2784
rect 2444 2696 2452 2704
rect 2428 2656 2436 2664
rect 2364 2636 2372 2644
rect 2412 2636 2420 2644
rect 2380 2616 2388 2624
rect 2348 2596 2356 2604
rect 2300 2556 2308 2564
rect 2332 2536 2340 2544
rect 2300 2496 2308 2504
rect 2332 2496 2340 2504
rect 2268 2396 2276 2404
rect 2284 2396 2292 2404
rect 2220 2336 2228 2344
rect 2236 2316 2244 2324
rect 2076 2296 2084 2304
rect 2092 2302 2100 2304
rect 2092 2296 2100 2302
rect 2156 2296 2164 2304
rect 2412 2576 2420 2584
rect 2540 3116 2548 3124
rect 2588 3116 2596 3124
rect 2700 3216 2708 3224
rect 2572 3076 2580 3084
rect 2540 3036 2548 3044
rect 2524 2996 2532 3004
rect 2508 2916 2516 2924
rect 2572 3036 2580 3044
rect 2620 3076 2628 3084
rect 2620 3036 2628 3044
rect 2636 3036 2644 3044
rect 2588 3016 2596 3024
rect 2604 3016 2612 3024
rect 2556 2996 2564 3004
rect 2684 3076 2692 3084
rect 2668 3036 2676 3044
rect 2652 3016 2660 3024
rect 2732 3176 2740 3184
rect 2828 3336 2836 3344
rect 2876 3356 2884 3364
rect 2876 3336 2884 3344
rect 2940 3416 2948 3424
rect 2956 3416 2964 3424
rect 2956 3396 2964 3404
rect 3020 3756 3028 3764
rect 3068 3816 3076 3824
rect 3113 3806 3121 3814
rect 3123 3806 3131 3814
rect 3133 3806 3141 3814
rect 3143 3806 3151 3814
rect 3084 3796 3092 3804
rect 3180 3796 3188 3804
rect 3260 4076 3268 4084
rect 3260 3896 3268 3904
rect 3260 3836 3268 3844
rect 3052 3756 3060 3764
rect 3004 3696 3012 3704
rect 3036 3696 3044 3704
rect 3068 3676 3076 3684
rect 3084 3676 3092 3684
rect 3132 3676 3140 3684
rect 3004 3656 3012 3664
rect 3068 3616 3076 3624
rect 3116 3616 3124 3624
rect 3068 3596 3076 3604
rect 3020 3556 3028 3564
rect 3036 3456 3044 3464
rect 3052 3436 3060 3444
rect 2988 3416 2996 3424
rect 2972 3376 2980 3384
rect 2940 3316 2948 3324
rect 2828 3256 2836 3264
rect 2844 3256 2852 3264
rect 2796 3236 2804 3244
rect 2780 3216 2788 3224
rect 2748 3136 2756 3144
rect 2780 3096 2788 3104
rect 2812 3216 2820 3224
rect 2796 3076 2804 3084
rect 2732 3056 2740 3064
rect 2748 2996 2756 3004
rect 2796 3036 2804 3044
rect 2812 2996 2820 3004
rect 2572 2936 2580 2944
rect 2508 2896 2516 2904
rect 2540 2896 2548 2904
rect 2556 2876 2564 2884
rect 2508 2856 2516 2864
rect 2508 2836 2516 2844
rect 2476 2776 2484 2784
rect 2492 2756 2500 2764
rect 2540 2776 2548 2784
rect 2588 2816 2596 2824
rect 2556 2736 2564 2744
rect 2572 2736 2580 2744
rect 2588 2736 2596 2744
rect 2764 2956 2772 2964
rect 2780 2956 2788 2964
rect 2636 2936 2644 2944
rect 2620 2896 2628 2904
rect 2604 2716 2612 2724
rect 2492 2696 2500 2704
rect 2524 2696 2532 2704
rect 2540 2696 2548 2704
rect 2684 2896 2692 2904
rect 2876 3236 2884 3244
rect 2860 3136 2868 3144
rect 2860 3116 2868 3124
rect 2988 3296 2996 3304
rect 3004 3296 3012 3304
rect 2892 3216 2900 3224
rect 2908 3216 2916 3224
rect 2940 3216 2948 3224
rect 2956 3216 2964 3224
rect 2972 3216 2980 3224
rect 2860 3076 2868 3084
rect 2876 3056 2884 3064
rect 2860 2996 2868 3004
rect 2748 2916 2756 2924
rect 2940 3136 2948 3144
rect 2972 3156 2980 3164
rect 2972 3116 2980 3124
rect 3004 3236 3012 3244
rect 3084 3576 3092 3584
rect 3100 3556 3108 3564
rect 3116 3456 3124 3464
rect 3148 3656 3156 3664
rect 3340 4136 3348 4144
rect 3356 4116 3364 4124
rect 3372 4076 3380 4084
rect 3596 4296 3604 4304
rect 3644 4296 3652 4304
rect 3420 4276 3428 4284
rect 3564 4276 3572 4284
rect 3580 4276 3588 4284
rect 3580 4256 3588 4264
rect 3420 4216 3428 4224
rect 3468 4216 3476 4224
rect 3436 4196 3444 4204
rect 3468 4116 3476 4124
rect 3564 4116 3572 4124
rect 3468 4076 3476 4084
rect 3564 4076 3572 4084
rect 3388 4056 3396 4064
rect 3548 3996 3556 4004
rect 3372 3916 3380 3924
rect 3420 3936 3428 3944
rect 3404 3916 3412 3924
rect 3452 3916 3460 3924
rect 3468 3916 3476 3924
rect 3404 3896 3412 3904
rect 3324 3836 3332 3844
rect 3324 3776 3332 3784
rect 3308 3756 3316 3764
rect 3260 3716 3268 3724
rect 3292 3716 3300 3724
rect 3308 3716 3316 3724
rect 3228 3696 3236 3704
rect 3260 3676 3268 3684
rect 3372 3756 3380 3764
rect 3388 3716 3396 3724
rect 3324 3656 3332 3664
rect 3340 3656 3348 3664
rect 3180 3596 3188 3604
rect 3324 3596 3332 3604
rect 3244 3556 3252 3564
rect 3308 3556 3316 3564
rect 3212 3536 3220 3544
rect 3228 3536 3236 3544
rect 3132 3436 3140 3444
rect 3292 3536 3300 3544
rect 3228 3436 3236 3444
rect 3084 3416 3092 3424
rect 3180 3416 3188 3424
rect 3113 3406 3121 3414
rect 3123 3406 3131 3414
rect 3133 3406 3141 3414
rect 3143 3406 3151 3414
rect 3180 3396 3188 3404
rect 3148 3376 3156 3384
rect 3084 3316 3092 3324
rect 3100 3296 3108 3304
rect 3036 3176 3044 3184
rect 3100 3176 3108 3184
rect 3052 3136 3060 3144
rect 3084 3096 3092 3104
rect 3180 3336 3188 3344
rect 3164 3316 3172 3324
rect 3260 3376 3268 3384
rect 3292 3376 3300 3384
rect 3148 3136 3156 3144
rect 3100 3076 3108 3084
rect 2972 3036 2980 3044
rect 2988 3036 2996 3044
rect 3068 3036 3076 3044
rect 3212 3296 3216 3304
rect 3216 3296 3220 3304
rect 3244 3296 3252 3304
rect 3212 3256 3220 3264
rect 3228 3256 3236 3264
rect 3196 3136 3204 3144
rect 3180 3076 3188 3084
rect 2908 3016 2916 3024
rect 2940 3016 2948 3024
rect 3004 2996 3012 3004
rect 2924 2956 2932 2964
rect 3068 2956 3076 2964
rect 2892 2936 2900 2944
rect 2908 2916 2916 2924
rect 2796 2836 2804 2844
rect 2748 2816 2756 2824
rect 2716 2776 2724 2784
rect 2652 2756 2660 2764
rect 2684 2756 2692 2764
rect 2700 2756 2708 2764
rect 2652 2716 2660 2724
rect 2460 2656 2468 2664
rect 2444 2556 2452 2564
rect 2508 2676 2516 2684
rect 2556 2656 2564 2664
rect 2508 2636 2516 2644
rect 2524 2636 2532 2644
rect 2396 2536 2404 2544
rect 2476 2536 2484 2544
rect 2492 2536 2500 2544
rect 2396 2496 2404 2504
rect 2428 2496 2436 2504
rect 2380 2476 2388 2484
rect 2412 2476 2420 2484
rect 2364 2436 2372 2444
rect 2396 2376 2404 2384
rect 2364 2356 2372 2364
rect 2364 2336 2372 2344
rect 2300 2316 2308 2324
rect 2172 2276 2180 2284
rect 2236 2276 2244 2284
rect 2316 2276 2324 2284
rect 2172 2256 2180 2264
rect 2268 2256 2276 2264
rect 2332 2256 2340 2264
rect 2156 2216 2164 2224
rect 2060 2196 2068 2204
rect 2108 2196 2116 2204
rect 2188 2196 2196 2204
rect 2268 2196 2276 2204
rect 2044 2176 2052 2184
rect 1996 2136 2004 2144
rect 2012 2136 2020 2144
rect 2012 2096 2020 2104
rect 1996 2076 2004 2084
rect 1980 1976 1988 1984
rect 2044 1976 2052 1984
rect 2012 1936 2020 1944
rect 1964 1896 1972 1904
rect 1980 1896 1988 1904
rect 1884 1856 1892 1864
rect 1900 1856 1908 1864
rect 1916 1856 1924 1864
rect 1868 1776 1876 1784
rect 1740 1656 1748 1664
rect 1708 1596 1716 1604
rect 1692 1576 1700 1584
rect 1676 1516 1684 1524
rect 1756 1596 1764 1604
rect 1756 1536 1764 1544
rect 1676 1496 1684 1504
rect 1740 1496 1748 1504
rect 1660 1456 1668 1464
rect 1724 1456 1732 1464
rect 1676 1436 1684 1444
rect 1612 1396 1620 1404
rect 1628 1396 1636 1404
rect 1740 1416 1748 1424
rect 1740 1396 1748 1404
rect 1612 1376 1620 1384
rect 1612 1356 1620 1364
rect 1660 1356 1668 1364
rect 1612 1336 1620 1344
rect 1644 1336 1652 1344
rect 1660 1316 1668 1324
rect 1596 1296 1604 1304
rect 1612 1296 1620 1304
rect 1644 1256 1652 1264
rect 1548 1216 1556 1224
rect 1577 1206 1585 1214
rect 1587 1206 1595 1214
rect 1597 1206 1605 1214
rect 1607 1206 1615 1214
rect 1548 1196 1556 1204
rect 1500 1136 1508 1144
rect 1516 1136 1524 1144
rect 1724 1176 1732 1184
rect 1708 1136 1716 1144
rect 1484 1116 1492 1124
rect 1532 1116 1540 1124
rect 1644 1116 1652 1124
rect 1772 1476 1780 1484
rect 1772 1456 1780 1464
rect 1804 1696 1812 1704
rect 1852 1736 1860 1744
rect 1980 1856 1988 1864
rect 2092 2156 2100 2164
rect 2060 1896 2068 1904
rect 2108 2096 2116 2104
rect 2156 2096 2164 2104
rect 2172 2096 2180 2104
rect 2172 2076 2180 2084
rect 2332 2156 2340 2164
rect 2204 2096 2212 2104
rect 2236 2096 2244 2104
rect 2412 2356 2420 2364
rect 2428 2336 2436 2344
rect 2428 2316 2436 2324
rect 2412 2196 2420 2204
rect 2220 1996 2228 2004
rect 2140 1976 2148 1984
rect 2172 1976 2180 1984
rect 2188 1976 2196 1984
rect 2332 2096 2340 2104
rect 2364 2036 2372 2044
rect 2332 2016 2340 2024
rect 2348 2016 2356 2024
rect 2380 2016 2388 2024
rect 2396 2016 2404 2024
rect 2124 1956 2132 1964
rect 1900 1736 1908 1744
rect 1884 1716 1892 1724
rect 1948 1836 1956 1844
rect 1980 1836 1988 1844
rect 1996 1836 2004 1844
rect 1932 1756 1940 1764
rect 2012 1816 2020 1824
rect 2044 1836 2052 1844
rect 2076 1836 2084 1844
rect 2028 1796 2036 1804
rect 2044 1796 2052 1804
rect 2060 1776 2068 1784
rect 2076 1776 2084 1784
rect 2044 1756 2052 1764
rect 1948 1736 1956 1744
rect 2028 1736 2036 1744
rect 1948 1716 1956 1724
rect 1916 1696 1924 1704
rect 1884 1656 1892 1664
rect 1932 1656 1940 1664
rect 1804 1536 1812 1544
rect 1820 1516 1828 1524
rect 1932 1596 1940 1604
rect 1980 1716 1988 1724
rect 1964 1676 1972 1684
rect 1964 1656 1972 1664
rect 2012 1696 2020 1704
rect 1980 1576 1988 1584
rect 1964 1516 1972 1524
rect 1900 1456 1908 1464
rect 1916 1456 1924 1464
rect 1948 1456 1956 1464
rect 1804 1416 1812 1424
rect 1900 1436 1908 1444
rect 1948 1436 1956 1444
rect 1884 1396 1892 1404
rect 1804 1356 1812 1364
rect 1852 1356 1860 1364
rect 1868 1356 1876 1364
rect 1788 1336 1796 1344
rect 1900 1356 1908 1364
rect 2044 1596 2052 1604
rect 2028 1576 2036 1584
rect 2012 1516 2020 1524
rect 2044 1496 2052 1504
rect 1820 1316 1828 1324
rect 1884 1316 1892 1324
rect 1804 1176 1812 1184
rect 1756 1116 1764 1124
rect 1676 1096 1684 1104
rect 1740 1096 1748 1104
rect 1788 1096 1796 1104
rect 1532 1076 1540 1084
rect 1612 1076 1620 1084
rect 1644 1076 1652 1084
rect 1388 996 1396 1004
rect 1420 996 1428 1004
rect 1372 976 1380 984
rect 1308 936 1316 944
rect 1292 876 1300 884
rect 1340 936 1348 944
rect 1516 1016 1524 1024
rect 1452 956 1460 964
rect 1468 956 1476 964
rect 1564 1056 1572 1064
rect 1564 1016 1572 1024
rect 1596 1016 1604 1024
rect 1580 956 1588 964
rect 1708 1076 1716 1084
rect 1804 1076 1812 1084
rect 1836 1276 1844 1284
rect 1852 1256 1860 1264
rect 1868 1196 1876 1204
rect 2028 1476 2036 1484
rect 2156 1936 2164 1944
rect 2220 1956 2228 1964
rect 2252 1956 2260 1964
rect 2172 1916 2180 1924
rect 2140 1896 2148 1904
rect 2236 1916 2244 1924
rect 2348 1976 2356 1984
rect 2332 1936 2340 1944
rect 2476 2376 2484 2384
rect 2460 2336 2468 2344
rect 2444 2256 2452 2264
rect 2652 2676 2660 2684
rect 2604 2656 2612 2664
rect 2636 2656 2644 2664
rect 2588 2556 2596 2564
rect 2636 2616 2644 2624
rect 2652 2616 2660 2624
rect 2620 2596 2628 2604
rect 2556 2536 2564 2544
rect 2604 2536 2612 2544
rect 2508 2376 2516 2384
rect 2492 2316 2500 2324
rect 2492 2276 2500 2284
rect 2460 2196 2468 2204
rect 2444 2176 2452 2184
rect 2492 2176 2500 2184
rect 2460 2156 2468 2164
rect 2476 2156 2484 2164
rect 2492 2156 2500 2164
rect 2556 2336 2564 2344
rect 2812 2756 2820 2764
rect 2796 2736 2804 2744
rect 2764 2716 2772 2724
rect 2684 2696 2692 2704
rect 2748 2696 2756 2704
rect 2684 2676 2692 2684
rect 2748 2676 2756 2684
rect 2684 2656 2692 2664
rect 2700 2636 2708 2644
rect 2748 2636 2756 2644
rect 2700 2596 2708 2604
rect 2636 2516 2644 2524
rect 2620 2496 2628 2504
rect 2604 2376 2612 2384
rect 2620 2376 2628 2384
rect 2588 2336 2596 2344
rect 2524 2316 2532 2324
rect 2572 2316 2580 2324
rect 2668 2376 2676 2384
rect 2636 2356 2644 2364
rect 2652 2356 2660 2364
rect 2796 2576 2804 2584
rect 2716 2556 2724 2564
rect 2764 2536 2772 2544
rect 2684 2336 2692 2344
rect 2588 2296 2596 2304
rect 2604 2296 2612 2304
rect 2540 2276 2548 2284
rect 2556 2276 2564 2284
rect 2524 2256 2532 2264
rect 2588 2276 2596 2284
rect 2652 2276 2660 2284
rect 2588 2256 2596 2264
rect 2668 2256 2676 2264
rect 2684 2256 2692 2264
rect 2556 2176 2564 2184
rect 2684 2176 2692 2184
rect 2604 2156 2612 2164
rect 2540 2096 2548 2104
rect 2572 2096 2580 2104
rect 2492 2016 2500 2024
rect 2540 2016 2548 2024
rect 2444 1976 2452 1984
rect 2476 1976 2484 1984
rect 2268 1876 2276 1884
rect 2284 1876 2292 1884
rect 2316 1876 2324 1884
rect 2204 1856 2212 1864
rect 2252 1856 2260 1864
rect 2140 1816 2148 1824
rect 2124 1736 2132 1744
rect 2092 1696 2100 1704
rect 2124 1696 2132 1704
rect 2092 1676 2100 1684
rect 2108 1656 2116 1664
rect 2092 1596 2100 1604
rect 2092 1576 2100 1584
rect 2060 1476 2068 1484
rect 2044 1456 2052 1464
rect 2108 1516 2116 1524
rect 2172 1816 2180 1824
rect 2188 1816 2196 1824
rect 2156 1796 2164 1804
rect 2156 1756 2164 1764
rect 2156 1576 2164 1584
rect 2172 1576 2180 1584
rect 2140 1536 2148 1544
rect 2140 1516 2148 1524
rect 2124 1476 2132 1484
rect 2140 1456 2148 1464
rect 2156 1456 2164 1464
rect 2028 1396 2036 1404
rect 2028 1356 2036 1364
rect 2028 1336 2036 1344
rect 2012 1316 2020 1324
rect 1948 1276 1956 1284
rect 1916 1256 1924 1264
rect 2028 1256 2036 1264
rect 1900 1236 1908 1244
rect 1884 1116 1892 1124
rect 2092 1396 2100 1404
rect 2108 1356 2116 1364
rect 2076 1316 2084 1324
rect 2092 1316 2100 1324
rect 2348 1876 2356 1884
rect 2364 1876 2372 1884
rect 2316 1816 2324 1824
rect 2380 1836 2388 1844
rect 2364 1796 2372 1804
rect 2428 1876 2436 1884
rect 2460 1876 2468 1884
rect 2476 1876 2484 1884
rect 2412 1836 2420 1844
rect 2380 1776 2388 1784
rect 2204 1736 2212 1744
rect 2220 1716 2228 1724
rect 2236 1716 2244 1724
rect 2204 1656 2212 1664
rect 2220 1656 2228 1664
rect 2220 1596 2228 1604
rect 2348 1756 2356 1764
rect 2300 1736 2308 1744
rect 2316 1716 2324 1724
rect 2268 1536 2276 1544
rect 2300 1596 2308 1604
rect 2460 1796 2468 1804
rect 2540 1976 2548 1984
rect 2604 2036 2612 2044
rect 2588 1956 2596 1964
rect 2540 1936 2548 1944
rect 2540 1916 2548 1924
rect 2716 2476 2724 2484
rect 2716 2396 2724 2404
rect 2780 2476 2788 2484
rect 2844 2716 2852 2724
rect 2844 2656 2852 2664
rect 2844 2556 2852 2564
rect 2892 2856 2900 2864
rect 2876 2836 2884 2844
rect 2892 2716 2900 2724
rect 2876 2616 2884 2624
rect 2876 2576 2884 2584
rect 2972 2936 2980 2944
rect 2940 2916 2948 2924
rect 2924 2756 2932 2764
rect 2940 2756 2948 2764
rect 2988 2916 2996 2924
rect 3036 2936 3044 2944
rect 3020 2916 3028 2924
rect 3052 2916 3060 2924
rect 3036 2876 3044 2884
rect 3068 2876 3076 2884
rect 2988 2856 2996 2864
rect 3020 2856 3028 2864
rect 2988 2836 2996 2844
rect 2924 2716 2932 2724
rect 2940 2716 2948 2724
rect 2972 2716 2980 2724
rect 2908 2696 2916 2704
rect 2908 2636 2916 2644
rect 3052 2856 3060 2864
rect 3164 3036 3172 3044
rect 3113 3006 3121 3014
rect 3123 3006 3131 3014
rect 3133 3006 3141 3014
rect 3143 3006 3151 3014
rect 3276 3316 3284 3324
rect 3260 3176 3268 3184
rect 3420 3716 3428 3724
rect 3404 3656 3412 3664
rect 3372 3616 3380 3624
rect 3388 3616 3396 3624
rect 3356 3556 3364 3564
rect 3388 3496 3396 3504
rect 3372 3456 3380 3464
rect 3372 3436 3380 3444
rect 3372 3356 3380 3364
rect 3420 3616 3428 3624
rect 3468 3876 3476 3884
rect 3484 3676 3492 3684
rect 3532 3936 3540 3944
rect 3644 4236 3652 4244
rect 3628 4196 3636 4204
rect 3644 4176 3652 4184
rect 3612 4136 3620 4144
rect 3964 4516 3972 4524
rect 4140 4516 4148 4524
rect 4252 4516 4260 4524
rect 4204 4496 4212 4504
rect 4140 4476 4148 4484
rect 3900 4456 3908 4464
rect 3948 4456 3956 4464
rect 3692 4356 3700 4364
rect 3772 4356 3780 4364
rect 3676 4336 3684 4344
rect 3884 4316 3892 4324
rect 3740 4196 3748 4204
rect 3996 4316 4004 4324
rect 4076 4316 4084 4324
rect 3788 4216 3796 4224
rect 3772 4196 3780 4204
rect 3996 4236 4004 4244
rect 3756 4176 3764 4184
rect 3964 4176 3972 4184
rect 3676 4156 3684 4164
rect 3724 4156 3732 4164
rect 3612 4116 3620 4124
rect 3660 4116 3668 4124
rect 3612 4096 3620 4104
rect 3596 4056 3604 4064
rect 3596 3996 3604 4004
rect 3612 3996 3620 4004
rect 3644 3996 3652 4004
rect 3580 3936 3588 3944
rect 3692 4136 3700 4144
rect 3820 4136 3828 4144
rect 3932 4136 3940 4144
rect 4092 4276 4100 4284
rect 4156 4276 4164 4284
rect 4124 4256 4132 4264
rect 4076 4216 4084 4224
rect 3708 4096 3716 4104
rect 3836 4096 3844 4104
rect 3916 4096 3924 4104
rect 3724 4076 3732 4084
rect 3852 4076 3860 4084
rect 3900 4076 3908 4084
rect 3900 3996 3908 4004
rect 4028 4136 4036 4144
rect 4044 4136 4052 4144
rect 4204 4296 4212 4304
rect 4204 4276 4212 4284
rect 4428 4496 4436 4504
rect 4540 4496 4548 4504
rect 4348 4456 4356 4464
rect 4508 4476 4516 4484
rect 4636 4516 4644 4524
rect 4732 4476 4740 4484
rect 4780 4476 4788 4484
rect 4540 4456 4548 4464
rect 4572 4456 4580 4464
rect 4860 4456 4868 4464
rect 4508 4416 4516 4424
rect 4284 4296 4292 4304
rect 4348 4296 4356 4304
rect 4444 4296 4452 4304
rect 4508 4296 4516 4304
rect 4268 4276 4276 4284
rect 4300 4276 4308 4284
rect 4188 4256 4196 4264
rect 4220 4256 4228 4264
rect 4252 4256 4260 4264
rect 4188 4236 4196 4244
rect 4172 4156 4180 4164
rect 4028 4116 4036 4124
rect 4092 4116 4100 4124
rect 4172 4096 4180 4104
rect 4076 4076 4084 4084
rect 4092 4076 4100 4084
rect 4044 3996 4052 4004
rect 4012 3956 4020 3964
rect 3948 3936 3956 3944
rect 3740 3916 3748 3924
rect 3548 3876 3556 3884
rect 3532 3776 3540 3784
rect 3516 3736 3524 3744
rect 3516 3716 3524 3724
rect 3452 3616 3460 3624
rect 3468 3556 3476 3564
rect 3532 3556 3540 3564
rect 3436 3496 3444 3504
rect 3452 3496 3460 3504
rect 3420 3456 3428 3464
rect 3420 3396 3428 3404
rect 3420 3336 3428 3344
rect 3228 3076 3236 3084
rect 3212 3036 3220 3044
rect 3228 3016 3236 3024
rect 3116 2956 3124 2964
rect 3180 2956 3188 2964
rect 3196 2956 3204 2964
rect 3100 2916 3108 2924
rect 3036 2816 3044 2824
rect 3004 2756 3012 2764
rect 3004 2736 3012 2744
rect 3084 2836 3092 2844
rect 3340 3316 3348 3324
rect 3404 3316 3412 3324
rect 3420 3316 3428 3324
rect 3356 3296 3364 3304
rect 3372 3296 3376 3304
rect 3376 3296 3380 3304
rect 3356 3236 3364 3244
rect 3340 3136 3348 3144
rect 3388 3236 3396 3244
rect 3388 3156 3396 3164
rect 3372 3116 3380 3124
rect 3388 3056 3396 3064
rect 3260 2996 3268 3004
rect 3340 3016 3348 3024
rect 3356 3016 3364 3024
rect 3308 2956 3316 2964
rect 3260 2936 3268 2944
rect 3324 2936 3332 2944
rect 3228 2916 3236 2924
rect 3180 2876 3188 2884
rect 3196 2876 3204 2884
rect 3116 2856 3124 2864
rect 3132 2856 3140 2864
rect 3244 2896 3252 2904
rect 3116 2836 3124 2844
rect 3068 2776 3076 2784
rect 3052 2736 3060 2744
rect 3068 2736 3076 2744
rect 3020 2716 3028 2724
rect 3100 2776 3108 2784
rect 2956 2596 2964 2604
rect 2828 2536 2836 2544
rect 2940 2536 2948 2544
rect 3116 2696 3124 2704
rect 3228 2836 3236 2844
rect 3164 2816 3172 2824
rect 3180 2796 3188 2804
rect 3164 2776 3172 2784
rect 3148 2716 3156 2724
rect 3212 2776 3220 2784
rect 3196 2736 3204 2744
rect 3004 2676 3012 2684
rect 3068 2676 3076 2684
rect 3100 2676 3108 2684
rect 3132 2676 3140 2684
rect 3180 2676 3188 2684
rect 2988 2616 2996 2624
rect 3100 2636 3108 2644
rect 3116 2636 3124 2644
rect 3052 2616 3060 2624
rect 3084 2616 3092 2624
rect 3180 2616 3188 2624
rect 3036 2596 3044 2604
rect 3068 2596 3076 2604
rect 2844 2496 2852 2504
rect 2860 2476 2868 2484
rect 2812 2436 2820 2444
rect 2828 2436 2836 2444
rect 2732 2376 2740 2384
rect 2828 2376 2836 2384
rect 2844 2376 2852 2384
rect 2796 2356 2804 2364
rect 2892 2496 2900 2504
rect 2876 2436 2884 2444
rect 2764 2316 2772 2324
rect 2780 2316 2788 2324
rect 2748 2296 2756 2304
rect 2748 2256 2756 2264
rect 2732 2216 2740 2224
rect 2876 2336 2884 2344
rect 2908 2476 2916 2484
rect 2924 2376 2932 2384
rect 2844 2276 2852 2284
rect 2876 2276 2884 2284
rect 2892 2276 2900 2284
rect 2908 2276 2916 2284
rect 2828 2256 2836 2264
rect 2796 2216 2804 2224
rect 2764 2196 2772 2204
rect 2716 2176 2724 2184
rect 2764 2176 2772 2184
rect 2796 2156 2804 2164
rect 2812 2156 2820 2164
rect 2748 2136 2756 2144
rect 2716 2096 2724 2104
rect 2732 2096 2740 2104
rect 2636 2036 2644 2044
rect 2620 2016 2628 2024
rect 2652 2016 2660 2024
rect 2716 2016 2724 2024
rect 2620 1996 2628 2004
rect 2716 1996 2724 2004
rect 2780 2096 2788 2104
rect 2796 2096 2804 2104
rect 2780 2076 2788 2084
rect 2812 2056 2820 2064
rect 2796 2016 2804 2024
rect 2812 2016 2820 2024
rect 2620 1916 2628 1924
rect 2636 1916 2644 1924
rect 2540 1836 2548 1844
rect 2556 1836 2564 1844
rect 2572 1796 2580 1804
rect 2588 1796 2596 1804
rect 2540 1756 2548 1764
rect 2588 1756 2596 1764
rect 2412 1736 2420 1744
rect 2508 1736 2516 1744
rect 2348 1596 2356 1604
rect 2364 1596 2372 1604
rect 2236 1516 2244 1524
rect 2332 1516 2340 1524
rect 2188 1476 2196 1484
rect 2412 1716 2420 1724
rect 2428 1716 2436 1724
rect 2444 1676 2452 1684
rect 2396 1656 2404 1664
rect 2412 1656 2420 1664
rect 2396 1516 2404 1524
rect 2476 1556 2484 1564
rect 2476 1536 2484 1544
rect 2268 1496 2276 1504
rect 2300 1496 2308 1504
rect 2364 1496 2372 1504
rect 2380 1496 2388 1504
rect 2460 1496 2468 1504
rect 2492 1496 2500 1504
rect 2508 1496 2516 1504
rect 2252 1476 2260 1484
rect 2284 1476 2292 1484
rect 2172 1396 2180 1404
rect 2188 1396 2196 1404
rect 2348 1476 2356 1484
rect 2332 1416 2340 1424
rect 2348 1416 2356 1424
rect 2300 1356 2308 1364
rect 2060 1276 2068 1284
rect 2060 1216 2068 1224
rect 2044 1176 2052 1184
rect 1852 1076 1860 1084
rect 1676 1036 1684 1044
rect 1676 1016 1684 1024
rect 1708 1016 1716 1024
rect 1644 976 1652 984
rect 1772 1056 1780 1064
rect 1788 1056 1796 1064
rect 1820 1056 1828 1064
rect 1740 1036 1748 1044
rect 1628 956 1636 964
rect 1676 956 1684 964
rect 1724 956 1732 964
rect 1532 916 1540 924
rect 1628 916 1636 924
rect 1388 896 1396 904
rect 1500 876 1508 884
rect 1516 876 1524 884
rect 1340 856 1348 864
rect 1372 856 1380 864
rect 1372 816 1380 824
rect 1276 736 1284 744
rect 1340 736 1348 744
rect 1388 796 1396 804
rect 1388 776 1396 784
rect 1468 796 1476 804
rect 1516 776 1524 784
rect 1548 876 1556 884
rect 1548 816 1556 824
rect 1577 806 1585 814
rect 1587 806 1595 814
rect 1597 806 1605 814
rect 1607 806 1615 814
rect 1836 1036 1844 1044
rect 1852 1036 1860 1044
rect 1756 996 1764 1004
rect 1772 996 1780 1004
rect 1772 956 1780 964
rect 1756 916 1764 924
rect 1388 756 1396 764
rect 1436 756 1444 764
rect 1292 696 1300 704
rect 972 656 980 664
rect 1036 676 1044 684
rect 1084 676 1092 684
rect 1116 676 1124 684
rect 1164 676 1172 684
rect 1260 676 1268 684
rect 1324 676 1332 684
rect 1372 676 1380 684
rect 956 616 964 624
rect 988 616 996 624
rect 1036 616 1044 624
rect 1100 636 1108 644
rect 988 576 996 584
rect 1052 576 1060 584
rect 908 556 916 564
rect 924 556 932 564
rect 956 556 964 564
rect 940 496 948 504
rect 956 496 964 504
rect 828 396 836 404
rect 876 396 884 404
rect 1084 416 1092 424
rect 1084 376 1092 384
rect 1052 336 1060 344
rect 1132 656 1140 664
rect 1164 656 1172 664
rect 1228 656 1236 664
rect 1116 596 1124 604
rect 1260 636 1268 644
rect 1276 616 1284 624
rect 1436 736 1444 744
rect 1468 736 1476 744
rect 1484 736 1492 744
rect 1532 756 1540 764
rect 1596 756 1604 764
rect 1644 756 1652 764
rect 1580 736 1588 744
rect 1468 676 1476 684
rect 1548 676 1556 684
rect 1196 576 1204 584
rect 1324 576 1332 584
rect 1388 576 1396 584
rect 1436 576 1444 584
rect 1148 536 1156 544
rect 1372 536 1380 544
rect 1404 536 1412 544
rect 1116 496 1124 504
rect 1148 496 1156 504
rect 1484 636 1492 644
rect 1532 636 1540 644
rect 1468 536 1476 544
rect 1484 536 1492 544
rect 1436 516 1444 524
rect 1452 516 1460 524
rect 1500 516 1508 524
rect 1164 416 1172 424
rect 1180 416 1188 424
rect 1148 376 1156 384
rect 1084 316 1092 324
rect 1100 316 1108 324
rect 812 296 820 304
rect 1148 296 1156 304
rect 1228 396 1236 404
rect 1228 376 1236 384
rect 1260 336 1268 344
rect 1180 316 1188 324
rect 1196 316 1204 324
rect 924 276 932 284
rect 1276 296 1284 304
rect 1212 276 1220 284
rect 892 256 900 264
rect 988 256 996 264
rect 876 216 884 224
rect 972 216 980 224
rect 860 156 868 164
rect 780 136 788 144
rect 300 116 308 124
rect 380 116 386 124
rect 386 116 388 124
rect 460 116 468 124
rect 924 176 932 184
rect 1052 196 1060 204
rect 924 136 932 144
rect 1004 136 1012 144
rect 1084 236 1092 244
rect 1116 236 1124 244
rect 1068 176 1076 184
rect 1084 156 1092 164
rect 844 116 852 124
rect 572 56 580 64
rect 828 96 836 104
rect 972 116 980 124
rect 1404 496 1412 504
rect 1484 496 1492 504
rect 1404 396 1412 404
rect 1420 396 1428 404
rect 1452 336 1460 344
rect 1404 316 1412 324
rect 1308 276 1316 284
rect 1324 276 1332 284
rect 1340 276 1348 284
rect 1308 256 1316 264
rect 1548 576 1556 584
rect 1644 736 1652 744
rect 1692 896 1700 904
rect 1708 896 1716 904
rect 1756 896 1764 904
rect 1676 796 1684 804
rect 1740 816 1748 824
rect 1692 736 1700 744
rect 1756 716 1764 724
rect 1756 696 1764 704
rect 1740 656 1748 664
rect 1820 1016 1828 1024
rect 1836 956 1844 964
rect 1836 916 1844 924
rect 1820 896 1828 904
rect 1916 1096 1924 1104
rect 1948 1096 1956 1104
rect 1964 1096 1972 1104
rect 1916 1036 1924 1044
rect 1900 1016 1908 1024
rect 1900 976 1908 984
rect 1964 1056 1972 1064
rect 2012 1096 2020 1104
rect 2060 1096 2068 1104
rect 2076 1076 2084 1084
rect 2012 1056 2020 1064
rect 2060 1056 2068 1064
rect 2076 1056 2084 1064
rect 1980 1016 1988 1024
rect 1996 1016 2004 1024
rect 1996 996 2004 1004
rect 1916 956 1924 964
rect 1948 956 1956 964
rect 1980 956 1988 964
rect 1884 896 1892 904
rect 1884 736 1892 744
rect 1660 636 1668 644
rect 1724 636 1732 644
rect 1756 636 1764 644
rect 1660 616 1668 624
rect 1660 576 1668 584
rect 1724 576 1732 584
rect 1628 556 1636 564
rect 1644 536 1652 544
rect 1532 516 1540 524
rect 1596 516 1604 524
rect 1612 456 1620 464
rect 1548 436 1556 444
rect 1580 436 1588 444
rect 1516 416 1524 424
rect 1516 336 1524 344
rect 1500 316 1508 324
rect 1577 406 1585 414
rect 1587 406 1595 414
rect 1597 406 1605 414
rect 1607 406 1615 414
rect 1692 536 1700 544
rect 1644 396 1652 404
rect 1580 356 1588 364
rect 1564 316 1572 324
rect 1532 296 1540 304
rect 1548 296 1556 304
rect 1404 280 1412 284
rect 1404 276 1412 280
rect 1500 276 1508 284
rect 1388 256 1396 264
rect 1436 256 1444 264
rect 1596 336 1604 344
rect 1644 336 1652 344
rect 1628 316 1636 324
rect 1660 316 1668 324
rect 1724 536 1732 544
rect 1740 536 1748 544
rect 1772 536 1780 544
rect 1852 716 1860 724
rect 1868 696 1876 704
rect 1852 616 1860 624
rect 1884 596 1892 604
rect 1932 856 1940 864
rect 1948 856 1956 864
rect 1996 916 2004 924
rect 2060 1016 2068 1024
rect 2044 976 2052 984
rect 1916 796 1924 804
rect 1948 756 1956 764
rect 2108 1236 2116 1244
rect 2124 1236 2132 1244
rect 2220 1336 2228 1344
rect 2316 1336 2324 1344
rect 2364 1396 2372 1404
rect 2156 1316 2164 1324
rect 2188 1316 2196 1324
rect 2140 1136 2148 1144
rect 2172 1296 2180 1304
rect 2172 1176 2180 1184
rect 2268 1236 2276 1244
rect 2220 1216 2228 1224
rect 2252 1216 2260 1224
rect 2124 1096 2132 1104
rect 2172 1116 2180 1124
rect 2092 1016 2100 1024
rect 2076 976 2084 984
rect 2060 956 2068 964
rect 2156 1076 2164 1084
rect 2156 1016 2164 1024
rect 2108 956 2116 964
rect 2124 956 2132 964
rect 2156 956 2164 964
rect 2220 1076 2228 1084
rect 2188 1056 2196 1064
rect 2204 1056 2212 1064
rect 2220 1056 2228 1064
rect 2188 1016 2196 1024
rect 2172 936 2180 944
rect 2092 916 2100 924
rect 2012 856 2020 864
rect 2044 856 2052 864
rect 2124 856 2132 864
rect 2044 816 2052 824
rect 1932 736 1940 744
rect 1996 736 2004 744
rect 2028 696 2036 704
rect 1868 536 1876 544
rect 1804 516 1812 524
rect 1900 536 1908 544
rect 1708 496 1716 504
rect 1836 496 1844 504
rect 1852 496 1860 504
rect 1740 396 1748 404
rect 1852 436 1860 444
rect 2060 736 2068 744
rect 2044 676 2052 684
rect 1948 656 1956 664
rect 1932 616 1940 624
rect 1964 616 1972 624
rect 2044 616 2052 624
rect 1964 596 1972 604
rect 1980 596 1988 604
rect 2172 916 2180 924
rect 2124 816 2132 824
rect 2140 816 2148 824
rect 2172 756 2180 764
rect 2300 1176 2308 1184
rect 2268 1076 2276 1084
rect 2316 1076 2324 1084
rect 2252 1056 2260 1064
rect 2268 1056 2276 1064
rect 2236 996 2244 1004
rect 2252 996 2260 1004
rect 2396 1376 2404 1384
rect 2380 1356 2388 1364
rect 2380 1316 2388 1324
rect 2364 1236 2372 1244
rect 2364 1216 2372 1224
rect 2380 1196 2388 1204
rect 2428 1456 2436 1464
rect 2492 1456 2500 1464
rect 2428 1416 2436 1424
rect 2444 1416 2452 1424
rect 2428 1316 2436 1324
rect 2524 1456 2532 1464
rect 2636 1876 2644 1884
rect 2748 1956 2756 1964
rect 2812 1976 2820 1984
rect 3052 2556 3060 2564
rect 3068 2556 3076 2564
rect 3113 2606 3121 2614
rect 3123 2606 3131 2614
rect 3133 2606 3141 2614
rect 3143 2606 3151 2614
rect 3196 2596 3204 2604
rect 3196 2576 3204 2584
rect 3180 2556 3188 2564
rect 2972 2436 2980 2444
rect 2988 2436 2996 2444
rect 2956 2416 2964 2424
rect 2940 2336 2948 2344
rect 3100 2496 3108 2504
rect 3084 2476 3092 2484
rect 3132 2476 3140 2484
rect 3036 2436 3044 2444
rect 3020 2416 3028 2424
rect 3004 2296 3012 2304
rect 2908 2256 2916 2264
rect 2924 2216 2932 2224
rect 2940 2216 2948 2224
rect 2972 2216 2980 2224
rect 2860 2176 2868 2184
rect 2876 2176 2884 2184
rect 2844 2156 2852 2164
rect 2876 2156 2884 2164
rect 3052 2356 3060 2364
rect 3036 2276 3044 2284
rect 3020 2256 3028 2264
rect 3004 2216 3012 2224
rect 2860 2076 2868 2084
rect 2860 2056 2868 2064
rect 2876 2056 2884 2064
rect 2844 1976 2852 1984
rect 2876 2016 2884 2024
rect 2892 2016 2900 2024
rect 2716 1876 2724 1884
rect 2732 1876 2740 1884
rect 2812 1876 2820 1884
rect 2700 1856 2708 1864
rect 2780 1856 2788 1864
rect 2812 1856 2820 1864
rect 2764 1836 2772 1844
rect 2812 1836 2820 1844
rect 2732 1816 2740 1824
rect 2716 1776 2724 1784
rect 2556 1716 2564 1724
rect 2604 1676 2612 1684
rect 2620 1676 2628 1684
rect 2588 1616 2596 1624
rect 2604 1616 2612 1624
rect 2588 1596 2596 1604
rect 2556 1556 2564 1564
rect 2588 1556 2596 1564
rect 2508 1416 2516 1424
rect 2492 1336 2500 1344
rect 2492 1296 2500 1304
rect 2444 1256 2452 1264
rect 2412 1236 2420 1244
rect 2444 1236 2452 1244
rect 2428 1196 2436 1204
rect 2364 1116 2372 1124
rect 2476 1216 2484 1224
rect 2460 1136 2468 1144
rect 2412 1116 2420 1124
rect 2444 1116 2452 1124
rect 2268 956 2276 964
rect 2204 916 2212 924
rect 2204 756 2212 764
rect 2204 736 2212 744
rect 2252 876 2260 884
rect 2236 756 2244 764
rect 2188 716 2196 724
rect 2092 696 2100 704
rect 2156 696 2164 704
rect 2172 696 2180 704
rect 2108 656 2116 664
rect 2108 636 2116 644
rect 2284 816 2292 824
rect 2284 796 2292 804
rect 2332 1036 2340 1044
rect 2380 1036 2388 1044
rect 2444 1076 2452 1084
rect 2460 1076 2468 1084
rect 2428 1056 2436 1064
rect 2396 1016 2404 1024
rect 2332 996 2340 1004
rect 2396 996 2404 1004
rect 2412 976 2420 984
rect 2588 1456 2596 1464
rect 2796 1776 2804 1784
rect 2764 1756 2772 1764
rect 2716 1696 2724 1704
rect 2700 1656 2708 1664
rect 2668 1616 2676 1624
rect 2684 1616 2692 1624
rect 2652 1556 2660 1564
rect 2636 1536 2644 1544
rect 2604 1416 2612 1424
rect 2556 1316 2564 1324
rect 2524 1296 2532 1304
rect 2508 1276 2516 1284
rect 2748 1656 2756 1664
rect 2716 1616 2724 1624
rect 2700 1556 2708 1564
rect 2652 1476 2660 1484
rect 2636 1376 2644 1384
rect 2716 1476 2724 1484
rect 2668 1416 2676 1424
rect 2700 1416 2708 1424
rect 2652 1356 2660 1364
rect 2652 1336 2660 1344
rect 2668 1336 2676 1344
rect 2684 1336 2692 1344
rect 2700 1336 2708 1344
rect 2620 1316 2628 1324
rect 2636 1316 2644 1324
rect 2588 1296 2596 1304
rect 2604 1296 2612 1304
rect 2588 1276 2596 1284
rect 2620 1276 2628 1284
rect 2652 1276 2660 1284
rect 2588 1236 2596 1244
rect 2540 1216 2548 1224
rect 2556 1216 2564 1224
rect 2508 1116 2516 1124
rect 2524 1116 2532 1124
rect 2588 1136 2596 1144
rect 2556 1116 2564 1124
rect 2652 1156 2660 1164
rect 2620 1136 2628 1144
rect 2492 1076 2500 1084
rect 2604 1096 2612 1104
rect 2716 1316 2724 1324
rect 2732 1176 2740 1184
rect 2700 1156 2708 1164
rect 2716 1156 2724 1164
rect 2780 1696 2788 1704
rect 2796 1696 2804 1704
rect 2860 1956 2868 1964
rect 2892 1956 2900 1964
rect 2956 2116 2964 2124
rect 2972 2116 2980 2124
rect 3100 2456 3108 2464
rect 3084 2336 3092 2344
rect 3276 2916 3284 2924
rect 3260 2836 3268 2844
rect 3244 2816 3252 2824
rect 3420 3256 3428 3264
rect 3596 3836 3604 3844
rect 3580 3736 3588 3744
rect 3612 3736 3620 3744
rect 3676 3896 3684 3904
rect 3692 3896 3700 3904
rect 3740 3896 3748 3904
rect 3756 3896 3764 3904
rect 3772 3796 3780 3804
rect 3676 3756 3684 3764
rect 3724 3756 3732 3764
rect 3612 3696 3620 3704
rect 3596 3636 3604 3644
rect 3612 3636 3620 3644
rect 3564 3556 3572 3564
rect 3452 3456 3460 3464
rect 3468 3436 3476 3444
rect 3484 3416 3492 3424
rect 3468 3376 3476 3384
rect 3452 3356 3460 3364
rect 3420 3236 3428 3244
rect 3436 3236 3444 3244
rect 3420 3156 3428 3164
rect 3468 3256 3476 3264
rect 3548 3456 3556 3464
rect 3660 3716 3668 3724
rect 3692 3516 3700 3524
rect 3740 3696 3748 3704
rect 3772 3756 3780 3764
rect 3788 3756 3796 3764
rect 3724 3556 3732 3564
rect 3660 3496 3668 3504
rect 3692 3496 3700 3504
rect 3708 3496 3716 3504
rect 3724 3496 3732 3504
rect 3628 3476 3636 3484
rect 3596 3416 3604 3424
rect 3516 3396 3524 3404
rect 3532 3356 3540 3364
rect 3548 3356 3556 3364
rect 3580 3356 3588 3364
rect 3612 3356 3620 3364
rect 3500 3336 3508 3344
rect 3548 3336 3556 3344
rect 3500 3316 3508 3324
rect 3484 3176 3492 3184
rect 3500 3176 3508 3184
rect 3420 3116 3428 3124
rect 3452 3116 3460 3124
rect 3484 3116 3492 3124
rect 3356 2956 3364 2964
rect 3388 2956 3396 2964
rect 3436 3056 3444 3064
rect 3468 3036 3476 3044
rect 3452 2976 3460 2984
rect 3468 2956 3476 2964
rect 3436 2936 3444 2944
rect 3436 2916 3444 2924
rect 3340 2876 3348 2884
rect 3372 2856 3380 2864
rect 3324 2836 3332 2844
rect 3356 2836 3364 2844
rect 3292 2776 3300 2784
rect 3308 2776 3316 2784
rect 3228 2716 3236 2724
rect 3260 2736 3268 2744
rect 3292 2736 3300 2744
rect 3292 2716 3300 2724
rect 3228 2576 3236 2584
rect 3388 2836 3396 2844
rect 3404 2836 3412 2844
rect 3356 2756 3364 2764
rect 3372 2756 3380 2764
rect 3452 2836 3460 2844
rect 3548 3196 3556 3204
rect 3676 3456 3684 3464
rect 3644 3436 3652 3444
rect 3660 3416 3668 3424
rect 3724 3456 3732 3464
rect 3756 3456 3764 3464
rect 3852 3836 3860 3844
rect 3804 3736 3812 3744
rect 3820 3736 3828 3744
rect 3820 3696 3828 3704
rect 3884 3796 3892 3804
rect 3852 3756 3860 3764
rect 3868 3736 3876 3744
rect 4012 3936 4020 3944
rect 4060 3936 4068 3944
rect 4156 3936 4164 3944
rect 4060 3916 4068 3924
rect 4124 3916 4132 3924
rect 3948 3856 3956 3864
rect 4060 3876 4068 3884
rect 4076 3876 4084 3884
rect 4092 3876 4100 3884
rect 3996 3836 4004 3844
rect 3980 3796 3988 3804
rect 3996 3796 4004 3804
rect 3964 3756 3972 3764
rect 4156 3856 4164 3864
rect 4284 4216 4292 4224
rect 4204 4116 4212 4124
rect 4236 4116 4244 4124
rect 4396 4196 4404 4204
rect 4396 4176 4404 4184
rect 4380 4156 4388 4164
rect 4316 4136 4324 4144
rect 4300 4116 4308 4124
rect 4665 4406 4673 4414
rect 4675 4406 4683 4414
rect 4685 4406 4693 4414
rect 4695 4406 4703 4414
rect 4556 4296 4564 4304
rect 4604 4296 4612 4304
rect 5100 4496 5108 4504
rect 5052 4456 5060 4464
rect 5020 4436 5028 4444
rect 5436 4536 5444 4544
rect 5532 4536 5540 4544
rect 5260 4518 5268 4524
rect 5260 4516 5268 4518
rect 5324 4516 5332 4524
rect 5324 4496 5332 4504
rect 5244 4456 5252 4464
rect 5148 4416 5156 4424
rect 5100 4316 5108 4324
rect 4700 4296 4708 4304
rect 4908 4296 4916 4304
rect 4956 4296 4964 4304
rect 5052 4296 5060 4304
rect 5068 4302 5076 4304
rect 5068 4296 5076 4302
rect 4684 4276 4692 4284
rect 4732 4276 4740 4284
rect 4748 4276 4756 4284
rect 4652 4256 4660 4264
rect 4620 4236 4628 4244
rect 4604 4216 4612 4224
rect 4860 4256 4868 4264
rect 5052 4176 5060 4184
rect 4716 4136 4724 4144
rect 4780 4136 4788 4144
rect 5084 4156 5092 4164
rect 5740 4536 5748 4544
rect 5884 4536 5892 4544
rect 5404 4516 5412 4524
rect 5548 4516 5556 4524
rect 5692 4516 5700 4524
rect 5756 4516 5764 4524
rect 5788 4516 5796 4524
rect 5420 4496 5428 4504
rect 5484 4496 5492 4504
rect 5612 4496 5620 4504
rect 5676 4496 5684 4504
rect 5756 4496 5764 4504
rect 5372 4376 5380 4384
rect 5228 4356 5236 4364
rect 5164 4316 5172 4324
rect 5452 4476 5460 4484
rect 5468 4356 5476 4364
rect 5404 4316 5412 4324
rect 5660 4476 5668 4484
rect 5500 4456 5508 4464
rect 5548 4456 5556 4464
rect 5580 4456 5588 4464
rect 5484 4336 5492 4344
rect 5180 4296 5188 4304
rect 5356 4296 5364 4304
rect 5516 4316 5524 4324
rect 5612 4436 5620 4444
rect 5628 4436 5636 4444
rect 5788 4456 5796 4464
rect 5740 4436 5748 4444
rect 5708 4356 5716 4364
rect 5756 4356 5764 4364
rect 5820 4356 5828 4364
rect 5788 4336 5796 4344
rect 5628 4316 5636 4324
rect 5164 4276 5172 4284
rect 5228 4276 5236 4284
rect 5372 4276 5380 4284
rect 5420 4276 5428 4284
rect 5580 4276 5588 4284
rect 5596 4276 5604 4284
rect 5116 4156 5124 4164
rect 4364 4116 4372 4124
rect 4588 4116 4596 4124
rect 4764 4116 4772 4124
rect 4956 4116 4964 4124
rect 5020 4116 5028 4124
rect 4332 4096 4340 4104
rect 4380 4096 4388 4104
rect 4220 3996 4228 4004
rect 4204 3936 4212 3944
rect 4236 3936 4244 3944
rect 4220 3916 4228 3924
rect 4268 4076 4276 4084
rect 4300 4076 4308 4084
rect 4284 3996 4292 4004
rect 4348 3996 4356 4004
rect 4284 3976 4292 3984
rect 4348 3976 4356 3984
rect 4268 3916 4276 3924
rect 4252 3896 4260 3904
rect 4348 3896 4356 3904
rect 4508 3896 4516 3904
rect 4284 3876 4292 3884
rect 4556 3876 4564 3884
rect 4188 3856 4196 3864
rect 4396 3836 4404 3844
rect 4156 3796 4164 3804
rect 4172 3796 4180 3804
rect 4188 3796 4196 3804
rect 4092 3756 4100 3764
rect 3948 3716 3956 3724
rect 3980 3716 3988 3724
rect 3836 3676 3844 3684
rect 3836 3596 3844 3604
rect 3820 3456 3828 3464
rect 3852 3456 3860 3464
rect 3772 3436 3780 3444
rect 3724 3416 3732 3424
rect 3740 3416 3748 3424
rect 3676 3396 3684 3404
rect 3692 3396 3700 3404
rect 3660 3356 3668 3364
rect 3644 3316 3652 3324
rect 3932 3616 3940 3624
rect 3916 3536 3924 3544
rect 3900 3516 3908 3524
rect 3916 3516 3924 3524
rect 3932 3496 3940 3504
rect 3772 3356 3780 3364
rect 3804 3356 3812 3364
rect 3820 3356 3828 3364
rect 3612 3116 3620 3124
rect 3692 3316 3700 3324
rect 4172 3736 4180 3744
rect 4140 3716 4148 3724
rect 4156 3716 4164 3724
rect 4060 3696 4068 3704
rect 4124 3696 4132 3704
rect 3980 3676 3988 3684
rect 4028 3596 4036 3604
rect 4060 3596 4068 3604
rect 3964 3556 3972 3564
rect 3980 3556 3988 3564
rect 3964 3516 3972 3524
rect 4060 3556 4068 3564
rect 4092 3556 4100 3564
rect 4252 3776 4260 3784
rect 4236 3736 4244 3744
rect 4220 3716 4228 3724
rect 4188 3676 4196 3684
rect 4748 4096 4756 4104
rect 4940 4096 4948 4104
rect 4700 4056 4708 4064
rect 4665 4006 4673 4014
rect 4675 4006 4683 4014
rect 4685 4006 4693 4014
rect 4695 4006 4703 4014
rect 4636 3996 4644 4004
rect 4764 3902 4772 3904
rect 5100 4116 5108 4124
rect 5052 3936 5060 3944
rect 5084 3936 5092 3944
rect 5244 4196 5252 4204
rect 5180 4176 5188 4184
rect 5340 4216 5348 4224
rect 5436 4256 5444 4264
rect 5660 4276 5668 4284
rect 6172 4576 6180 4584
rect 5932 4556 5940 4564
rect 5996 4556 6004 4564
rect 6012 4556 6020 4564
rect 6060 4556 6068 4564
rect 6092 4556 6100 4564
rect 5932 4516 5940 4524
rect 5884 4416 5892 4424
rect 5868 4376 5876 4384
rect 5980 4476 5988 4484
rect 6156 4536 6164 4544
rect 6012 4476 6020 4484
rect 6108 4496 6116 4504
rect 6172 4496 6180 4504
rect 6060 4436 6068 4444
rect 6044 4416 6052 4424
rect 5996 4396 6004 4404
rect 6028 4396 6036 4404
rect 6076 4376 6084 4384
rect 5916 4356 5924 4364
rect 5948 4356 5956 4364
rect 6028 4356 6036 4364
rect 5852 4336 5860 4344
rect 5868 4336 5876 4344
rect 5884 4336 5892 4344
rect 5916 4336 5924 4344
rect 5756 4276 5764 4284
rect 5612 4256 5620 4264
rect 5692 4256 5700 4264
rect 5724 4256 5732 4264
rect 5740 4256 5748 4264
rect 5788 4256 5796 4264
rect 5388 4216 5396 4224
rect 5276 4176 5284 4184
rect 5388 4176 5396 4184
rect 5244 4136 5252 4144
rect 5260 4136 5268 4144
rect 5468 4156 5476 4164
rect 5500 4216 5508 4224
rect 5548 4176 5556 4184
rect 5660 4176 5668 4184
rect 5404 4136 5412 4144
rect 5900 4316 5908 4324
rect 5932 4296 5940 4304
rect 5900 4276 5908 4284
rect 5852 4236 5860 4244
rect 5804 4216 5812 4224
rect 5852 4196 5860 4204
rect 5564 4136 5572 4144
rect 5692 4136 5700 4144
rect 5740 4136 5748 4144
rect 5788 4136 5796 4144
rect 5244 4116 5252 4124
rect 5324 4116 5332 4124
rect 5372 4116 5380 4124
rect 5436 4116 5444 4124
rect 5484 4116 5492 4124
rect 5148 4096 5156 4104
rect 5228 4096 5236 4104
rect 5292 4096 5300 4104
rect 5324 4096 5332 4104
rect 5356 4096 5364 4104
rect 5212 4056 5220 4064
rect 5180 4016 5188 4024
rect 4988 3916 4996 3924
rect 5068 3916 5076 3924
rect 5196 3916 5204 3924
rect 4764 3896 4772 3902
rect 4796 3876 4804 3884
rect 4940 3876 4948 3884
rect 4588 3816 4596 3824
rect 4620 3816 4628 3824
rect 4700 3816 4708 3824
rect 4556 3756 4564 3764
rect 4300 3736 4308 3744
rect 4556 3736 4564 3744
rect 4284 3716 4292 3724
rect 4460 3716 4468 3724
rect 4252 3676 4260 3684
rect 4236 3556 4244 3564
rect 4252 3556 4260 3564
rect 4204 3536 4212 3544
rect 4108 3516 4116 3524
rect 3948 3436 3956 3444
rect 3964 3436 3972 3444
rect 3980 3416 3988 3424
rect 4236 3516 4244 3524
rect 4380 3616 4388 3624
rect 4380 3556 4388 3564
rect 4316 3516 4324 3524
rect 4220 3496 4228 3504
rect 4044 3436 4052 3444
rect 4124 3436 4132 3444
rect 4172 3436 4180 3444
rect 4268 3436 4276 3444
rect 4060 3336 4068 3344
rect 4076 3336 4084 3344
rect 4108 3336 4116 3344
rect 3884 3316 3892 3324
rect 3756 3236 3764 3244
rect 3772 3236 3780 3244
rect 3740 3196 3748 3204
rect 3660 3156 3668 3164
rect 3676 3156 3684 3164
rect 3692 3156 3700 3164
rect 3708 3116 3716 3124
rect 3532 3076 3540 3084
rect 3580 3076 3588 3084
rect 3644 3056 3652 3064
rect 3580 3036 3588 3044
rect 3596 2956 3604 2964
rect 3612 2936 3620 2944
rect 3500 2916 3508 2924
rect 3692 3076 3700 3084
rect 3820 3296 3828 3304
rect 3932 3276 3940 3284
rect 3804 3236 3812 3244
rect 3772 3136 3780 3144
rect 3788 3136 3796 3144
rect 3820 3136 3828 3144
rect 3772 3076 3780 3084
rect 3852 3196 3860 3204
rect 3868 3196 3876 3204
rect 3852 3136 3860 3144
rect 3884 3116 3892 3124
rect 4028 3296 4036 3304
rect 3964 3236 3972 3244
rect 4092 3236 4100 3244
rect 4092 3156 4100 3164
rect 4268 3416 4276 3424
rect 4140 3396 4148 3404
rect 4204 3396 4212 3404
rect 4156 3336 4164 3344
rect 4236 3336 4244 3344
rect 4172 3316 4180 3324
rect 4124 3196 4132 3204
rect 4140 3196 4148 3204
rect 4540 3716 4548 3724
rect 4604 3716 4612 3724
rect 4588 3696 4596 3704
rect 4588 3596 4596 3604
rect 4972 3816 4980 3824
rect 4908 3756 4916 3764
rect 4636 3736 4644 3744
rect 4876 3736 4884 3744
rect 5052 3896 5060 3904
rect 5052 3876 5060 3884
rect 5100 3876 5108 3884
rect 5116 3876 5124 3884
rect 5084 3796 5092 3804
rect 5164 3896 5172 3904
rect 5420 4056 5428 4064
rect 5484 4056 5492 4064
rect 5372 3996 5380 4004
rect 5244 3916 5252 3924
rect 5324 3916 5332 3924
rect 5340 3896 5348 3904
rect 5404 3916 5412 3924
rect 5436 3916 5444 3924
rect 5452 3896 5460 3904
rect 5468 3896 5476 3904
rect 5548 4116 5556 4124
rect 5772 4116 5780 4124
rect 5676 4096 5684 4104
rect 5756 4016 5764 4024
rect 5740 3936 5748 3944
rect 5196 3876 5204 3884
rect 5228 3876 5236 3884
rect 5244 3876 5252 3884
rect 5292 3876 5300 3884
rect 5404 3876 5412 3884
rect 5596 3896 5604 3904
rect 5676 3916 5684 3924
rect 5660 3896 5668 3904
rect 5708 3896 5716 3904
rect 5180 3856 5188 3864
rect 5244 3856 5252 3864
rect 5532 3856 5540 3864
rect 5628 3856 5636 3864
rect 5356 3836 5364 3844
rect 5260 3816 5268 3824
rect 5132 3796 5140 3804
rect 5196 3796 5204 3804
rect 5276 3796 5284 3804
rect 5244 3756 5252 3764
rect 4940 3736 4948 3744
rect 5036 3716 5044 3724
rect 5148 3716 5156 3724
rect 4828 3696 4836 3704
rect 4636 3616 4644 3624
rect 4665 3606 4673 3614
rect 4675 3606 4683 3614
rect 4685 3606 4693 3614
rect 4695 3606 4703 3614
rect 4588 3556 4596 3564
rect 4556 3516 4564 3524
rect 4588 3516 4596 3524
rect 4732 3536 4740 3544
rect 4732 3516 4740 3524
rect 4892 3516 4900 3524
rect 4556 3496 4564 3504
rect 4460 3436 4468 3444
rect 4300 3376 4308 3384
rect 4332 3376 4340 3384
rect 4796 3496 4804 3504
rect 4844 3496 4852 3504
rect 4860 3496 4868 3504
rect 4780 3456 4788 3464
rect 4348 3336 4356 3344
rect 4476 3336 4484 3344
rect 4604 3336 4612 3344
rect 4748 3376 4756 3384
rect 4764 3376 4772 3384
rect 4732 3336 4740 3344
rect 4268 3316 4276 3324
rect 4316 3316 4324 3324
rect 4316 3296 4324 3304
rect 4412 3296 4420 3304
rect 4428 3296 4436 3304
rect 4236 3216 4244 3224
rect 3980 3136 3988 3144
rect 3996 3136 4004 3144
rect 4028 3136 4036 3144
rect 4172 3136 4180 3144
rect 4636 3276 4644 3284
rect 4476 3256 4484 3264
rect 4108 3116 4116 3124
rect 4124 3116 4132 3124
rect 4156 3116 4164 3124
rect 4188 3116 4192 3124
rect 4192 3116 4196 3124
rect 3948 3096 3956 3104
rect 4044 3096 4052 3104
rect 3868 3076 3876 3084
rect 3660 2996 3668 3004
rect 3692 2996 3700 3004
rect 3756 2996 3764 3004
rect 3676 2956 3684 2964
rect 3724 2956 3732 2964
rect 3692 2936 3700 2944
rect 3548 2896 3556 2904
rect 3596 2896 3604 2904
rect 3612 2896 3620 2904
rect 3644 2896 3652 2904
rect 3660 2896 3668 2904
rect 3708 2896 3716 2904
rect 3548 2856 3556 2864
rect 3580 2816 3588 2824
rect 3516 2796 3524 2804
rect 3564 2796 3572 2804
rect 3612 2836 3620 2844
rect 3660 2836 3668 2844
rect 3436 2736 3444 2744
rect 3452 2716 3460 2724
rect 3308 2656 3316 2664
rect 3356 2656 3364 2664
rect 3276 2636 3284 2644
rect 3292 2636 3300 2644
rect 3260 2576 3268 2584
rect 3244 2556 3252 2564
rect 3228 2476 3236 2484
rect 3212 2456 3220 2464
rect 3180 2396 3188 2404
rect 3196 2396 3204 2404
rect 3116 2316 3124 2324
rect 3100 2296 3108 2304
rect 3116 2296 3124 2304
rect 3116 2256 3124 2264
rect 3228 2416 3236 2424
rect 3228 2376 3236 2384
rect 3228 2256 3236 2264
rect 3100 2236 3108 2244
rect 3212 2236 3220 2244
rect 3084 2216 3092 2224
rect 3212 2216 3220 2224
rect 3068 2156 3076 2164
rect 2988 2096 2996 2104
rect 3004 2096 3012 2104
rect 2940 2076 2948 2084
rect 3020 2076 3028 2084
rect 2988 2056 2996 2064
rect 2972 2016 2980 2024
rect 2940 1936 2948 1944
rect 2924 1896 2932 1904
rect 2956 1876 2964 1884
rect 2876 1796 2884 1804
rect 3036 2056 3044 2064
rect 3113 2206 3121 2214
rect 3123 2206 3131 2214
rect 3133 2206 3141 2214
rect 3143 2206 3151 2214
rect 3180 2196 3188 2204
rect 3100 2176 3108 2184
rect 3084 2136 3092 2144
rect 3100 1976 3108 1984
rect 3100 1956 3108 1964
rect 3228 2136 3236 2144
rect 3132 2096 3140 2104
rect 3148 2096 3156 2104
rect 3164 2076 3172 2084
rect 3180 2016 3188 2024
rect 3196 2016 3204 2024
rect 3100 1916 3108 1924
rect 3116 1916 3124 1924
rect 3036 1896 3044 1904
rect 3084 1896 3092 1904
rect 2972 1836 2980 1844
rect 3180 1976 3188 1984
rect 3212 1976 3220 1984
rect 3180 1856 3188 1864
rect 3113 1806 3121 1814
rect 3123 1806 3131 1814
rect 3133 1806 3141 1814
rect 3143 1806 3151 1814
rect 2844 1776 2852 1784
rect 3084 1776 3092 1784
rect 2972 1756 2980 1764
rect 2988 1756 2996 1764
rect 2828 1736 2836 1744
rect 2860 1736 2868 1744
rect 2940 1736 2948 1744
rect 2876 1716 2884 1724
rect 2812 1676 2820 1684
rect 2860 1696 2868 1704
rect 2844 1676 2852 1684
rect 2892 1656 2900 1664
rect 2908 1656 2916 1664
rect 2828 1616 2836 1624
rect 2860 1616 2868 1624
rect 2860 1596 2868 1604
rect 2764 1516 2772 1524
rect 2796 1516 2804 1524
rect 2780 1496 2788 1504
rect 2812 1496 2820 1504
rect 2844 1516 2852 1524
rect 2828 1476 2836 1484
rect 2764 1416 2772 1424
rect 2780 1376 2788 1384
rect 2828 1356 2836 1364
rect 2892 1476 2900 1484
rect 2892 1436 2900 1444
rect 2876 1416 2884 1424
rect 2860 1376 2868 1384
rect 2796 1336 2804 1344
rect 2812 1336 2820 1344
rect 2844 1336 2852 1344
rect 2780 1316 2788 1324
rect 2876 1316 2884 1324
rect 2476 1056 2484 1064
rect 2540 1056 2548 1064
rect 2460 1036 2468 1044
rect 2476 1036 2484 1044
rect 2620 1036 2628 1044
rect 2348 956 2356 964
rect 2412 956 2420 964
rect 2428 956 2436 964
rect 2316 876 2324 884
rect 2300 756 2308 764
rect 2332 816 2340 824
rect 2172 676 2180 684
rect 2156 656 2164 664
rect 2172 636 2180 644
rect 2188 636 2196 644
rect 2236 676 2244 684
rect 2268 656 2276 664
rect 2108 596 2116 604
rect 2124 596 2132 604
rect 1996 556 2004 564
rect 2076 556 2084 564
rect 1916 496 1924 504
rect 1948 496 1956 504
rect 1884 436 1892 444
rect 1868 396 1876 404
rect 1884 396 1892 404
rect 1612 276 1620 284
rect 1692 296 1700 304
rect 1724 316 1732 324
rect 1884 316 1892 324
rect 1900 316 1908 324
rect 1708 276 1716 284
rect 1740 276 1748 284
rect 1868 296 1876 304
rect 1932 456 1940 464
rect 1980 456 1988 464
rect 2012 456 2020 464
rect 2044 456 2052 464
rect 2060 456 2068 464
rect 2124 576 2132 584
rect 2236 596 2244 604
rect 2156 556 2164 564
rect 2188 556 2196 564
rect 2172 536 2180 544
rect 2204 536 2212 544
rect 2140 496 2148 504
rect 2156 496 2164 504
rect 2188 516 2196 524
rect 2252 536 2260 544
rect 2332 656 2340 664
rect 2380 856 2388 864
rect 2396 836 2404 844
rect 2428 856 2436 864
rect 2668 996 2676 1004
rect 2540 956 2548 964
rect 2556 956 2564 964
rect 2588 956 2596 964
rect 2652 956 2660 964
rect 2476 836 2484 844
rect 2524 896 2532 904
rect 2588 896 2596 904
rect 2556 856 2564 864
rect 2540 776 2548 784
rect 2476 756 2484 764
rect 2492 756 2500 764
rect 2444 736 2452 744
rect 2460 736 2468 744
rect 2460 696 2468 704
rect 2524 736 2532 744
rect 2396 676 2404 684
rect 2444 676 2452 684
rect 2364 576 2372 584
rect 2364 556 2372 564
rect 2380 556 2388 564
rect 2316 536 2324 544
rect 2284 516 2292 524
rect 2300 516 2308 524
rect 2220 496 2228 504
rect 2444 576 2452 584
rect 2572 736 2580 744
rect 2604 736 2612 744
rect 2588 716 2596 724
rect 2556 656 2564 664
rect 2524 636 2532 644
rect 2540 636 2548 644
rect 2380 536 2388 544
rect 2348 516 2356 524
rect 2364 516 2372 524
rect 2428 516 2436 524
rect 2204 456 2212 464
rect 2220 456 2228 464
rect 2332 456 2340 464
rect 2140 436 2148 444
rect 2140 416 2148 424
rect 2236 416 2244 424
rect 2252 416 2260 424
rect 1932 296 1940 304
rect 2028 296 2036 304
rect 2092 296 2100 304
rect 1724 256 1732 264
rect 1356 236 1364 244
rect 1548 236 1556 244
rect 1580 236 1588 244
rect 1596 236 1604 244
rect 1196 196 1204 204
rect 1244 196 1252 204
rect 1276 196 1284 204
rect 1292 196 1300 204
rect 1340 196 1348 204
rect 1164 176 1172 184
rect 1180 176 1188 184
rect 1292 156 1300 164
rect 1516 196 1524 204
rect 1388 156 1396 164
rect 1484 156 1492 164
rect 1164 136 1172 144
rect 1292 136 1300 144
rect 1324 136 1332 144
rect 1372 136 1380 144
rect 1244 116 1252 124
rect 1276 116 1284 124
rect 1356 116 1364 124
rect 908 96 916 104
rect 1068 96 1076 104
rect 1132 96 1140 104
rect 1228 96 1236 104
rect 1308 96 1316 104
rect 876 76 884 84
rect 1020 76 1028 84
rect 1052 76 1060 84
rect 1660 216 1668 224
rect 1692 216 1700 224
rect 1708 216 1716 224
rect 1708 176 1716 184
rect 1724 176 1732 184
rect 1452 116 1460 124
rect 1500 116 1508 124
rect 1564 116 1572 124
rect 1580 116 1588 124
rect 1404 96 1412 104
rect 1420 96 1428 104
rect 1452 76 1460 84
rect 1580 76 1588 84
rect 1596 76 1604 84
rect 1644 116 1652 124
rect 1660 116 1668 124
rect 1788 276 1796 284
rect 1884 276 1892 284
rect 1900 276 1908 284
rect 1932 276 1940 284
rect 1996 256 2004 264
rect 2188 336 2196 344
rect 2236 336 2244 344
rect 2156 316 2164 324
rect 2236 316 2244 324
rect 2188 296 2196 304
rect 2316 416 2324 424
rect 2476 536 2484 544
rect 2492 496 2500 504
rect 2460 436 2468 444
rect 2396 396 2404 404
rect 2332 336 2340 344
rect 2332 296 2340 304
rect 2364 316 2372 324
rect 2460 356 2468 364
rect 2492 316 2500 324
rect 2364 296 2372 304
rect 2524 536 2532 544
rect 2060 256 2068 264
rect 2076 256 2084 264
rect 2012 236 2020 244
rect 1884 216 1892 224
rect 1836 196 1844 204
rect 1916 216 1924 224
rect 1932 216 1940 224
rect 1964 216 1972 224
rect 1980 216 1988 224
rect 1804 116 1812 124
rect 1900 116 1908 124
rect 1852 96 1860 104
rect 1932 96 1940 104
rect 1948 96 1956 104
rect 1980 176 1988 184
rect 2044 196 2052 204
rect 2060 176 2068 184
rect 2060 156 2068 164
rect 2028 116 2036 124
rect 2124 236 2132 244
rect 2204 236 2212 244
rect 2252 236 2260 244
rect 2156 196 2164 204
rect 2172 196 2180 204
rect 2092 156 2100 164
rect 2108 156 2116 164
rect 2204 156 2212 164
rect 2252 156 2260 164
rect 2076 116 2084 124
rect 1996 96 2004 104
rect 2028 76 2036 84
rect 2092 96 2100 104
rect 2140 136 2148 144
rect 2156 136 2164 144
rect 2220 136 2228 144
rect 2572 636 2580 644
rect 2556 616 2564 624
rect 2572 616 2580 624
rect 2588 616 2596 624
rect 2588 596 2596 604
rect 2620 596 2628 604
rect 2604 576 2612 584
rect 2620 556 2628 564
rect 2652 836 2660 844
rect 2748 1116 2756 1124
rect 2780 1276 2788 1284
rect 2732 1076 2740 1084
rect 2748 1076 2756 1084
rect 2764 1036 2772 1044
rect 2812 1276 2820 1284
rect 2860 1276 2868 1284
rect 2796 1196 2804 1204
rect 2812 1196 2820 1204
rect 2796 1036 2804 1044
rect 2828 1136 2836 1144
rect 2812 956 2820 964
rect 2716 776 2724 784
rect 2684 696 2692 704
rect 2652 676 2660 684
rect 2700 676 2708 684
rect 2668 656 2676 664
rect 2700 616 2708 624
rect 2780 796 2788 804
rect 2764 756 2772 764
rect 2780 676 2788 684
rect 2764 656 2772 664
rect 2812 796 2820 804
rect 2860 956 2868 964
rect 2924 1616 2932 1624
rect 2924 1596 2932 1604
rect 3212 1856 3220 1864
rect 3212 1836 3220 1844
rect 3260 2276 3268 2284
rect 3244 2076 3252 2084
rect 3308 2576 3316 2584
rect 3564 2756 3572 2764
rect 3596 2756 3604 2764
rect 3516 2716 3524 2724
rect 3532 2716 3540 2724
rect 3548 2716 3556 2724
rect 3468 2656 3476 2664
rect 3452 2616 3460 2624
rect 3404 2596 3412 2604
rect 3532 2636 3540 2644
rect 3500 2616 3508 2624
rect 3516 2616 3524 2624
rect 3468 2596 3476 2604
rect 3484 2596 3492 2604
rect 3324 2556 3332 2564
rect 3372 2556 3380 2564
rect 3452 2556 3460 2564
rect 3292 2536 3300 2544
rect 3324 2536 3332 2544
rect 3372 2536 3380 2544
rect 3324 2396 3332 2404
rect 3292 2376 3300 2384
rect 3372 2456 3380 2464
rect 3484 2576 3492 2584
rect 3500 2576 3508 2584
rect 3500 2536 3508 2544
rect 3468 2476 3476 2484
rect 3484 2476 3492 2484
rect 3388 2436 3396 2444
rect 3420 2436 3428 2444
rect 3452 2436 3460 2444
rect 3340 2336 3348 2344
rect 3388 2336 3396 2344
rect 3308 2236 3316 2244
rect 3340 2236 3348 2244
rect 3372 2216 3380 2224
rect 3596 2716 3604 2724
rect 3836 3036 3844 3044
rect 3868 3036 3876 3044
rect 3932 3076 3940 3084
rect 3900 2976 3908 2984
rect 3932 2976 3940 2984
rect 3788 2916 3796 2924
rect 3804 2856 3812 2864
rect 3964 2936 3972 2944
rect 3980 2916 3988 2924
rect 4012 2916 4020 2924
rect 3868 2856 3876 2864
rect 3916 2896 3924 2904
rect 3948 2896 3956 2904
rect 4012 2896 4020 2904
rect 4012 2876 4020 2884
rect 3772 2796 3780 2804
rect 3836 2796 3844 2804
rect 3852 2796 3860 2804
rect 3884 2796 3892 2804
rect 3900 2796 3908 2804
rect 3724 2776 3732 2784
rect 3772 2776 3780 2784
rect 3740 2756 3748 2764
rect 3756 2756 3764 2764
rect 3724 2696 3732 2704
rect 3948 2756 3956 2764
rect 3852 2716 3860 2724
rect 4076 3076 4084 3084
rect 4076 2976 4084 2984
rect 4092 2976 4100 2984
rect 4060 2936 4068 2944
rect 4092 2916 4100 2924
rect 4124 2916 4132 2924
rect 4060 2856 4068 2864
rect 4044 2776 4052 2784
rect 4044 2736 4052 2744
rect 3788 2696 3796 2704
rect 3804 2696 3812 2704
rect 4044 2696 4052 2704
rect 3676 2656 3684 2664
rect 3692 2656 3700 2664
rect 3612 2636 3620 2644
rect 3564 2596 3572 2604
rect 3564 2576 3572 2584
rect 3772 2676 3780 2684
rect 3804 2676 3812 2684
rect 3756 2656 3764 2664
rect 3660 2596 3668 2604
rect 3724 2596 3732 2604
rect 3580 2536 3588 2544
rect 3564 2476 3572 2484
rect 3532 2436 3540 2444
rect 3580 2436 3588 2444
rect 3628 2436 3636 2444
rect 3564 2376 3572 2384
rect 3612 2376 3620 2384
rect 3836 2676 3844 2684
rect 3916 2676 3924 2684
rect 4012 2676 4020 2684
rect 4028 2676 4036 2684
rect 3868 2656 3876 2664
rect 3916 2656 3924 2664
rect 4012 2656 4020 2664
rect 3804 2596 3812 2604
rect 3820 2596 3828 2604
rect 3852 2596 3860 2604
rect 3692 2556 3700 2564
rect 3804 2556 3812 2564
rect 3836 2556 3844 2564
rect 3692 2496 3700 2504
rect 3996 2616 4004 2624
rect 3996 2576 4004 2584
rect 3996 2556 4004 2564
rect 3932 2536 3940 2544
rect 3868 2516 3876 2524
rect 3916 2516 3924 2524
rect 3836 2496 3844 2504
rect 3756 2476 3764 2484
rect 3788 2476 3796 2484
rect 3676 2436 3684 2444
rect 3660 2416 3668 2424
rect 3740 2416 3748 2424
rect 3644 2356 3652 2364
rect 3516 2280 3524 2284
rect 3516 2276 3524 2280
rect 3532 2276 3540 2284
rect 3468 2256 3476 2264
rect 3548 2256 3556 2264
rect 3420 2236 3428 2244
rect 3452 2236 3460 2244
rect 3484 2236 3492 2244
rect 3516 2236 3524 2244
rect 3388 2176 3396 2184
rect 3372 2156 3380 2164
rect 3468 2216 3476 2224
rect 3516 2176 3524 2184
rect 3564 2176 3572 2184
rect 3484 2156 3492 2164
rect 3420 2136 3428 2144
rect 3516 2136 3524 2144
rect 3532 2136 3540 2144
rect 3612 2296 3620 2304
rect 3628 2276 3636 2284
rect 3596 2256 3604 2264
rect 3644 2256 3652 2264
rect 3692 2256 3700 2264
rect 3724 2256 3732 2264
rect 3660 2236 3668 2244
rect 3724 2236 3732 2244
rect 3740 2236 3748 2244
rect 3916 2496 3924 2504
rect 3884 2476 3892 2484
rect 3964 2516 3972 2524
rect 3948 2496 3956 2504
rect 3868 2456 3876 2464
rect 3852 2436 3860 2444
rect 3932 2436 3940 2444
rect 3980 2436 3988 2444
rect 4012 2516 4020 2524
rect 4076 2756 4084 2764
rect 4076 2736 4084 2744
rect 4060 2556 4068 2564
rect 4028 2436 4036 2444
rect 3916 2396 3924 2404
rect 3996 2396 4004 2404
rect 4028 2396 4036 2404
rect 3836 2376 3844 2384
rect 3900 2376 3908 2384
rect 3868 2316 3876 2324
rect 3884 2276 3892 2284
rect 3916 2336 3924 2344
rect 4300 3096 4308 3104
rect 4348 3096 4356 3104
rect 4220 3076 4228 3084
rect 4268 3076 4276 3084
rect 4332 3076 4340 3084
rect 4204 3016 4212 3024
rect 4284 3016 4292 3024
rect 4284 2976 4292 2984
rect 4172 2936 4180 2944
rect 4268 2936 4276 2944
rect 4156 2796 4164 2804
rect 4236 2776 4244 2784
rect 4284 2776 4292 2784
rect 4284 2756 4292 2764
rect 4108 2656 4116 2664
rect 4236 2616 4244 2624
rect 4236 2596 4244 2604
rect 4172 2576 4180 2584
rect 4204 2576 4212 2584
rect 4140 2536 4148 2544
rect 4268 2696 4276 2704
rect 4284 2556 4292 2564
rect 4092 2516 4100 2524
rect 4108 2516 4116 2524
rect 4108 2496 4116 2504
rect 4092 2436 4100 2444
rect 3932 2296 3940 2304
rect 4060 2296 4068 2304
rect 3996 2276 4004 2284
rect 3820 2256 3828 2264
rect 3852 2256 3860 2264
rect 3900 2256 3908 2264
rect 3692 2216 3700 2224
rect 3612 2176 3620 2184
rect 3644 2156 3652 2164
rect 3500 2116 3508 2124
rect 3564 2116 3572 2124
rect 3324 2096 3332 2104
rect 3356 2096 3364 2104
rect 3260 2016 3268 2024
rect 3292 2016 3300 2024
rect 3276 1996 3284 2004
rect 3260 1936 3268 1944
rect 3244 1916 3252 1924
rect 3356 2056 3364 2064
rect 3340 1976 3348 1984
rect 3372 1996 3380 2004
rect 3356 1936 3364 1944
rect 3340 1916 3348 1924
rect 3260 1876 3268 1884
rect 3276 1876 3284 1884
rect 3276 1856 3284 1864
rect 3196 1776 3204 1784
rect 3244 1816 3252 1824
rect 3260 1816 3268 1824
rect 3212 1756 3220 1764
rect 3308 1836 3316 1844
rect 3292 1816 3300 1824
rect 3292 1796 3300 1804
rect 3356 1896 3364 1904
rect 3340 1876 3348 1884
rect 3628 2116 3636 2124
rect 3692 2116 3700 2124
rect 3612 2096 3620 2104
rect 3676 2096 3684 2104
rect 3724 2116 3732 2124
rect 3548 1996 3556 2004
rect 3580 1996 3588 2004
rect 3596 1996 3604 2004
rect 3420 1936 3428 1944
rect 3388 1916 3396 1924
rect 3388 1896 3396 1904
rect 3388 1876 3396 1884
rect 3404 1876 3412 1884
rect 3372 1856 3380 1864
rect 3324 1816 3332 1824
rect 3372 1816 3380 1824
rect 3324 1796 3332 1804
rect 3356 1796 3364 1804
rect 3388 1796 3396 1804
rect 3628 2016 3636 2024
rect 3612 1956 3620 1964
rect 3516 1916 3524 1924
rect 3532 1916 3540 1924
rect 3436 1896 3444 1904
rect 3516 1896 3524 1904
rect 3564 1896 3572 1904
rect 3596 1896 3604 1904
rect 3548 1876 3556 1884
rect 3596 1856 3604 1864
rect 3468 1816 3476 1824
rect 3420 1796 3428 1804
rect 3436 1796 3444 1804
rect 3356 1756 3364 1764
rect 3388 1756 3396 1764
rect 3420 1756 3428 1764
rect 3372 1716 3380 1724
rect 3388 1716 3396 1724
rect 3212 1676 3220 1684
rect 3228 1676 3236 1684
rect 3260 1676 3268 1684
rect 3100 1536 3108 1544
rect 3116 1536 3124 1544
rect 3244 1536 3252 1544
rect 3260 1536 3268 1544
rect 2972 1516 2980 1524
rect 3132 1516 3140 1524
rect 2940 1476 2948 1484
rect 2988 1456 2996 1464
rect 3004 1456 3012 1464
rect 3036 1456 3044 1464
rect 2940 1436 2948 1444
rect 2908 1376 2916 1384
rect 2892 1036 2900 1044
rect 2860 936 2868 944
rect 3004 1416 3012 1424
rect 2972 1376 2980 1384
rect 2988 1376 2996 1384
rect 2988 1356 2996 1364
rect 3100 1496 3108 1504
rect 3196 1476 3204 1484
rect 3100 1456 3108 1464
rect 3164 1456 3172 1464
rect 3068 1396 3076 1404
rect 3113 1406 3121 1414
rect 3123 1406 3131 1414
rect 3133 1406 3141 1414
rect 3143 1406 3151 1414
rect 3228 1456 3236 1464
rect 3196 1436 3204 1444
rect 3180 1396 3188 1404
rect 3260 1476 3268 1484
rect 3308 1476 3316 1484
rect 3132 1376 3140 1384
rect 3148 1376 3156 1384
rect 3084 1356 3092 1364
rect 3116 1356 3124 1364
rect 2972 1316 2980 1324
rect 3020 1276 3028 1284
rect 3036 1276 3044 1284
rect 2940 1216 2948 1224
rect 2972 1216 2980 1224
rect 2940 1116 2948 1124
rect 2924 1036 2932 1044
rect 2908 936 2916 944
rect 2924 916 2932 924
rect 2860 896 2868 904
rect 3084 1176 3092 1184
rect 3068 1156 3076 1164
rect 3020 1136 3028 1144
rect 3052 1136 3060 1144
rect 2956 1056 2964 1064
rect 3084 1136 3092 1144
rect 3164 1336 3172 1344
rect 3244 1316 3252 1324
rect 3180 1296 3188 1304
rect 3164 1276 3172 1284
rect 3180 1276 3188 1284
rect 3148 1196 3156 1204
rect 3164 1196 3172 1204
rect 3132 1176 3140 1184
rect 3212 1196 3220 1204
rect 3196 1176 3204 1184
rect 3084 1076 3092 1084
rect 3100 1076 3108 1084
rect 2972 1016 2980 1024
rect 2972 956 2980 964
rect 3020 1016 3028 1024
rect 3036 976 3044 984
rect 3004 936 3012 944
rect 2988 916 2996 924
rect 2988 896 2996 904
rect 2844 856 2852 864
rect 2908 856 2916 864
rect 2924 856 2932 864
rect 2940 856 2948 864
rect 2972 856 2980 864
rect 3020 876 3028 884
rect 3068 1036 3076 1044
rect 3084 1016 3092 1024
rect 3113 1006 3121 1014
rect 3123 1006 3131 1014
rect 3133 1006 3141 1014
rect 3143 1006 3151 1014
rect 3084 996 3092 1004
rect 3068 956 3076 964
rect 3100 956 3108 964
rect 3132 956 3140 964
rect 3052 936 3060 944
rect 3084 936 3092 944
rect 3068 916 3076 924
rect 3068 896 3076 904
rect 3084 876 3092 884
rect 3100 876 3108 884
rect 3052 856 3060 864
rect 2940 816 2948 824
rect 2844 796 2852 804
rect 2828 736 2836 744
rect 2828 716 2836 724
rect 2908 716 2912 724
rect 2912 716 2916 724
rect 2812 656 2820 664
rect 2780 636 2788 644
rect 2796 636 2804 644
rect 3100 836 3108 844
rect 3116 836 3124 844
rect 3020 796 3028 804
rect 3068 796 3076 804
rect 3084 796 3092 804
rect 3004 736 3012 744
rect 2924 696 2932 704
rect 2972 696 2980 704
rect 2860 616 2868 624
rect 2972 656 2980 664
rect 2972 636 2980 644
rect 2892 616 2900 624
rect 2876 596 2884 604
rect 2844 576 2852 584
rect 2860 556 2868 564
rect 2636 536 2644 544
rect 2748 536 2756 544
rect 2780 536 2788 544
rect 2828 536 2836 544
rect 2572 516 2580 524
rect 2588 516 2596 524
rect 2636 516 2644 524
rect 2748 516 2756 524
rect 2572 496 2580 504
rect 2988 536 2996 544
rect 2908 516 2916 524
rect 2972 516 2980 524
rect 2652 496 2660 504
rect 2812 496 2820 504
rect 2844 496 2852 504
rect 2556 436 2564 444
rect 2604 436 2612 444
rect 2540 336 2548 344
rect 2540 316 2548 324
rect 2572 336 2580 344
rect 2620 336 2628 344
rect 2636 336 2644 344
rect 2668 336 2676 344
rect 2604 316 2612 324
rect 2668 316 2676 324
rect 2620 296 2628 304
rect 2524 256 2532 264
rect 2396 216 2404 224
rect 2412 216 2420 224
rect 2652 276 2660 284
rect 2556 216 2564 224
rect 2572 216 2580 224
rect 2716 356 2724 364
rect 2748 416 2756 424
rect 2924 496 2932 504
rect 3068 676 3076 684
rect 3020 616 3028 624
rect 3340 1456 3348 1464
rect 3452 1576 3460 1584
rect 3436 1536 3444 1544
rect 3580 1776 3588 1784
rect 3500 1756 3508 1764
rect 3564 1756 3572 1764
rect 3500 1716 3508 1724
rect 3468 1556 3476 1564
rect 3452 1476 3460 1484
rect 3452 1456 3460 1464
rect 3388 1416 3396 1424
rect 3292 1396 3300 1404
rect 3372 1396 3380 1404
rect 3468 1436 3476 1444
rect 3436 1396 3444 1404
rect 3452 1396 3460 1404
rect 3420 1376 3428 1384
rect 3388 1336 3396 1344
rect 3276 1316 3284 1324
rect 3292 1316 3300 1324
rect 3340 1296 3348 1304
rect 3292 1256 3300 1264
rect 3292 1136 3300 1144
rect 3308 1136 3316 1144
rect 3260 1116 3268 1124
rect 3244 1076 3252 1084
rect 3292 1076 3300 1084
rect 3292 1056 3300 1064
rect 3244 996 3252 1004
rect 3276 956 3284 964
rect 3372 1276 3380 1284
rect 3420 1296 3428 1304
rect 3388 1256 3396 1264
rect 3372 1096 3380 1104
rect 3500 1536 3508 1544
rect 3660 1996 3668 2004
rect 3676 1996 3684 2004
rect 3756 2216 3764 2224
rect 3756 2136 3764 2144
rect 3884 2196 3892 2204
rect 3820 2156 3828 2164
rect 3836 2156 3844 2164
rect 3788 2116 3796 2124
rect 3772 2096 3780 2104
rect 3804 1996 3812 2004
rect 3676 1936 3684 1944
rect 3708 1936 3716 1944
rect 3740 1936 3748 1944
rect 3644 1916 3652 1924
rect 3788 1916 3796 1924
rect 3660 1856 3668 1864
rect 3724 1856 3732 1864
rect 3740 1856 3748 1864
rect 3612 1756 3620 1764
rect 3660 1796 3668 1804
rect 3532 1596 3540 1604
rect 3580 1596 3588 1604
rect 3612 1596 3620 1604
rect 3628 1596 3636 1604
rect 3548 1576 3556 1584
rect 3564 1576 3572 1584
rect 3564 1496 3572 1504
rect 3628 1496 3636 1504
rect 3644 1476 3652 1484
rect 3564 1456 3572 1464
rect 3628 1456 3636 1464
rect 3516 1436 3524 1444
rect 3500 1316 3508 1324
rect 3532 1318 3540 1324
rect 3532 1316 3540 1318
rect 3484 1276 3492 1284
rect 3532 1276 3540 1284
rect 3516 1116 3524 1124
rect 3420 1076 3428 1084
rect 3404 1016 3412 1024
rect 3372 976 3380 984
rect 3388 976 3396 984
rect 3388 956 3396 964
rect 3212 936 3220 944
rect 3340 936 3348 944
rect 3196 916 3204 924
rect 3228 896 3236 904
rect 3196 876 3204 884
rect 3244 836 3252 844
rect 3340 896 3348 904
rect 3308 736 3316 744
rect 3244 716 3252 724
rect 3260 716 3268 724
rect 3308 716 3316 724
rect 3196 696 3204 704
rect 3212 696 3220 704
rect 3132 676 3140 684
rect 3084 656 3092 664
rect 3100 656 3108 664
rect 3148 656 3156 664
rect 3068 556 3076 564
rect 3113 606 3121 614
rect 3123 606 3131 614
rect 3133 606 3141 614
rect 3143 606 3151 614
rect 3180 596 3188 604
rect 3116 576 3124 584
rect 3164 576 3172 584
rect 3132 556 3140 564
rect 3100 536 3108 544
rect 3020 516 3028 524
rect 3036 516 3044 524
rect 3084 516 3092 524
rect 3116 516 3124 524
rect 3068 496 3076 504
rect 2908 396 2916 404
rect 2972 396 2980 404
rect 2732 336 2740 344
rect 2828 336 2836 344
rect 2876 336 2884 344
rect 2764 316 2772 324
rect 2748 296 2756 304
rect 2700 276 2708 284
rect 2716 276 2724 284
rect 2828 316 2836 324
rect 2940 336 2948 344
rect 2972 336 2980 344
rect 2924 316 2932 324
rect 2956 316 2964 324
rect 2988 316 2996 324
rect 2908 296 2916 304
rect 2908 276 2916 284
rect 2924 276 2932 284
rect 2972 276 2980 284
rect 3292 696 3300 704
rect 3228 636 3236 644
rect 3228 616 3236 624
rect 3228 576 3236 584
rect 3260 616 3268 624
rect 3228 556 3236 564
rect 3244 556 3252 564
rect 3292 556 3300 564
rect 3420 976 3428 984
rect 3404 876 3412 884
rect 3628 1376 3636 1384
rect 3564 1216 3572 1224
rect 3564 1196 3572 1204
rect 3532 1096 3540 1104
rect 3516 1076 3524 1084
rect 3596 1236 3604 1244
rect 3612 1156 3620 1164
rect 3580 1096 3588 1104
rect 3484 1036 3492 1044
rect 3468 1016 3476 1024
rect 3484 1016 3492 1024
rect 3548 1036 3556 1044
rect 3516 996 3524 1004
rect 3756 1796 3764 1804
rect 3676 1756 3684 1764
rect 3692 1756 3700 1764
rect 3868 2136 3876 2144
rect 3900 2176 3908 2184
rect 3852 2116 3860 2124
rect 3868 2116 3876 2124
rect 3820 1976 3828 1984
rect 3852 1936 3860 1944
rect 3804 1876 3812 1884
rect 3820 1876 3828 1884
rect 3772 1756 3780 1764
rect 3804 1756 3812 1764
rect 3916 2156 3924 2164
rect 3932 2136 3940 2144
rect 3932 2096 3940 2104
rect 3964 2096 3972 2104
rect 3980 2096 3988 2104
rect 4060 2096 4068 2104
rect 4076 2096 4084 2104
rect 3996 2056 4004 2064
rect 4012 2056 4020 2064
rect 3964 1976 3972 1984
rect 3996 1976 4004 1984
rect 3980 1916 3988 1924
rect 4028 2036 4036 2044
rect 4044 1996 4052 2004
rect 4044 1956 4052 1964
rect 4060 1956 4068 1964
rect 4044 1916 4052 1924
rect 4012 1876 4020 1884
rect 4060 1876 4068 1884
rect 3900 1816 3908 1824
rect 3836 1796 3844 1804
rect 3852 1796 3860 1804
rect 3900 1756 3908 1764
rect 4028 1836 4036 1844
rect 3980 1756 3988 1764
rect 4012 1756 4020 1764
rect 3740 1716 3748 1724
rect 3724 1556 3732 1564
rect 3708 1496 3716 1504
rect 3820 1716 3828 1724
rect 3932 1736 3940 1744
rect 3932 1696 3940 1704
rect 3964 1696 3972 1704
rect 4012 1676 4020 1684
rect 4012 1616 4020 1624
rect 3900 1556 3908 1564
rect 3932 1516 3940 1524
rect 3980 1516 3988 1524
rect 3916 1496 3924 1504
rect 3948 1496 3956 1504
rect 4012 1496 4020 1504
rect 4044 1816 4052 1824
rect 4044 1616 4052 1624
rect 4140 2496 4148 2504
rect 4172 2496 4180 2504
rect 4252 2496 4260 2504
rect 4428 3096 4436 3104
rect 4412 3076 4420 3084
rect 4460 3076 4468 3084
rect 4508 3196 4516 3204
rect 4524 3096 4532 3104
rect 4396 3036 4404 3044
rect 4428 3036 4436 3044
rect 4460 3036 4468 3044
rect 4508 3036 4516 3044
rect 4348 3016 4356 3024
rect 4316 2936 4324 2944
rect 4492 3016 4500 3024
rect 4380 2956 4388 2964
rect 4572 2956 4580 2964
rect 4540 2936 4548 2944
rect 4348 2916 4356 2924
rect 4348 2696 4356 2704
rect 4316 2656 4324 2664
rect 4300 2516 4308 2524
rect 4236 2436 4244 2444
rect 4268 2436 4276 2444
rect 4124 2376 4132 2384
rect 4156 2336 4164 2344
rect 4188 2336 4196 2344
rect 4124 2316 4132 2324
rect 4204 2296 4212 2304
rect 4284 2416 4292 2424
rect 4300 2416 4308 2424
rect 4396 2916 4404 2924
rect 4524 2916 4532 2924
rect 4665 3206 4673 3214
rect 4675 3206 4683 3214
rect 4685 3206 4693 3214
rect 4695 3206 4703 3214
rect 4668 3136 4676 3144
rect 4892 3376 4900 3384
rect 4780 3316 4788 3324
rect 4796 3316 4804 3324
rect 4844 3316 4852 3324
rect 4860 3316 4868 3324
rect 4844 3296 4852 3304
rect 4892 3296 4900 3304
rect 4796 3136 4804 3144
rect 4780 3116 4788 3124
rect 4844 3116 4852 3124
rect 4876 3096 4884 3104
rect 4700 3076 4708 3084
rect 4732 3076 4740 3084
rect 4732 3036 4740 3044
rect 4652 2976 4660 2984
rect 4652 2956 4660 2964
rect 4636 2936 4644 2944
rect 4636 2916 4644 2924
rect 4396 2736 4404 2744
rect 4684 2936 4692 2944
rect 4732 2936 4740 2944
rect 4860 2916 4868 2924
rect 5004 3696 5012 3704
rect 5116 3696 5124 3704
rect 5148 3696 5156 3704
rect 5180 3736 5188 3744
rect 5228 3716 5236 3724
rect 5084 3636 5092 3644
rect 5164 3636 5172 3644
rect 5180 3636 5188 3644
rect 4956 3496 4964 3504
rect 5228 3616 5236 3624
rect 5196 3576 5204 3584
rect 5420 3816 5428 3824
rect 5372 3756 5380 3764
rect 5388 3736 5396 3744
rect 5372 3716 5380 3724
rect 5356 3696 5364 3704
rect 5372 3696 5380 3704
rect 5324 3616 5332 3624
rect 5356 3616 5364 3624
rect 5308 3596 5316 3604
rect 5452 3796 5460 3804
rect 5676 3816 5684 3824
rect 5740 3796 5748 3804
rect 5660 3776 5668 3784
rect 5436 3756 5444 3764
rect 5516 3756 5524 3764
rect 5724 3756 5732 3764
rect 5452 3736 5460 3744
rect 5468 3736 5476 3744
rect 5436 3716 5444 3724
rect 5468 3676 5476 3684
rect 5452 3636 5460 3644
rect 5276 3576 5284 3584
rect 5324 3576 5332 3584
rect 5420 3576 5428 3584
rect 5244 3536 5252 3544
rect 5116 3516 5124 3524
rect 5084 3476 5092 3484
rect 5132 3476 5140 3484
rect 5180 3476 5188 3484
rect 5116 3416 5124 3424
rect 5308 3536 5316 3544
rect 5244 3476 5252 3484
rect 5260 3476 5268 3484
rect 5276 3456 5284 3464
rect 5276 3436 5284 3444
rect 5228 3396 5236 3404
rect 5292 3396 5300 3404
rect 5244 3356 5252 3364
rect 5292 3356 5300 3364
rect 4956 3336 4964 3344
rect 5004 3316 5012 3324
rect 5004 3096 5012 3104
rect 5180 3336 5188 3344
rect 5228 3336 5236 3344
rect 5052 3316 5060 3324
rect 5116 3316 5124 3324
rect 5164 3316 5172 3324
rect 5372 3516 5380 3524
rect 5836 4116 5844 4124
rect 5788 3996 5796 4004
rect 5788 3956 5796 3964
rect 5772 3936 5780 3944
rect 5932 4276 5940 4284
rect 5948 4256 5956 4264
rect 5916 4236 5924 4244
rect 5980 4236 5988 4244
rect 5996 4216 6004 4224
rect 5916 4196 5924 4204
rect 5948 4196 5956 4204
rect 6044 4256 6052 4264
rect 5980 4156 5988 4164
rect 5884 4116 5892 4124
rect 5900 4116 5908 4124
rect 5852 4016 5860 4024
rect 5916 4096 5924 4104
rect 6028 4196 6036 4204
rect 6092 4256 6100 4264
rect 6060 4176 6068 4184
rect 6060 4156 6068 4164
rect 6140 4436 6148 4444
rect 6124 4336 6132 4344
rect 6156 4416 6164 4424
rect 6204 4496 6212 4504
rect 6188 4436 6196 4444
rect 6284 4456 6292 4464
rect 6236 4416 6244 4424
rect 6172 4356 6180 4364
rect 6204 4356 6212 4364
rect 6124 4176 6132 4184
rect 6044 4136 6052 4144
rect 6028 4116 6036 4124
rect 5932 4076 5940 4084
rect 5980 4036 5988 4044
rect 5852 3996 5860 4004
rect 5884 3996 5892 4004
rect 5948 4016 5956 4024
rect 5964 3996 5972 4004
rect 5900 3976 5908 3984
rect 5932 3956 5940 3964
rect 5884 3936 5892 3944
rect 5900 3936 5908 3944
rect 5836 3916 5844 3924
rect 5820 3896 5828 3904
rect 5868 3896 5876 3904
rect 5772 3876 5780 3884
rect 5836 3876 5844 3884
rect 5916 3896 5924 3904
rect 5948 3916 5956 3924
rect 5836 3856 5844 3864
rect 5868 3856 5876 3864
rect 5788 3836 5796 3844
rect 5804 3796 5812 3804
rect 5516 3716 5524 3724
rect 5532 3716 5540 3724
rect 5580 3716 5588 3724
rect 5628 3716 5636 3724
rect 5724 3716 5732 3724
rect 5724 3696 5732 3704
rect 5756 3696 5764 3704
rect 5484 3656 5492 3664
rect 5548 3656 5556 3664
rect 5516 3636 5524 3644
rect 5676 3676 5684 3684
rect 5724 3676 5732 3684
rect 5788 3716 5796 3724
rect 5756 3656 5764 3664
rect 5772 3656 5780 3664
rect 5500 3616 5508 3624
rect 5564 3616 5572 3624
rect 5580 3616 5588 3624
rect 5596 3616 5604 3624
rect 5548 3556 5556 3564
rect 5500 3536 5508 3544
rect 5468 3496 5476 3504
rect 5532 3496 5540 3504
rect 5564 3516 5572 3524
rect 5788 3596 5796 3604
rect 5772 3516 5780 3524
rect 5580 3496 5588 3504
rect 5628 3496 5636 3504
rect 5676 3496 5684 3504
rect 5484 3476 5492 3484
rect 5644 3476 5652 3484
rect 5660 3476 5668 3484
rect 5340 3456 5348 3464
rect 5404 3456 5412 3464
rect 5420 3436 5428 3444
rect 5324 3416 5332 3424
rect 5452 3396 5460 3404
rect 5436 3376 5444 3384
rect 5516 3376 5524 3384
rect 5388 3356 5396 3364
rect 5324 3316 5332 3324
rect 5340 3316 5348 3324
rect 5084 3296 5092 3304
rect 5116 3296 5124 3304
rect 5196 3296 5204 3304
rect 5244 3296 5252 3304
rect 5340 3296 5348 3304
rect 5356 3296 5364 3304
rect 5420 3316 5428 3324
rect 5100 3236 5108 3244
rect 5388 3236 5396 3244
rect 5084 3156 5092 3164
rect 5052 3096 5060 3104
rect 4972 2956 4980 2964
rect 4908 2936 4916 2944
rect 5036 2936 5044 2944
rect 5020 2916 5028 2924
rect 4892 2876 4900 2884
rect 5020 2876 5028 2884
rect 4620 2836 4628 2844
rect 4636 2836 4644 2844
rect 4684 2836 4692 2844
rect 4620 2756 4628 2764
rect 4476 2696 4484 2704
rect 4492 2696 4500 2704
rect 4396 2656 4404 2664
rect 4444 2656 4452 2664
rect 4364 2576 4372 2584
rect 4364 2516 4372 2524
rect 4332 2436 4340 2444
rect 4252 2376 4260 2384
rect 4284 2376 4292 2384
rect 4156 2276 4164 2284
rect 4236 2276 4244 2284
rect 4140 2256 4148 2264
rect 4284 2256 4292 2264
rect 4284 2236 4292 2244
rect 4252 2176 4260 2184
rect 4124 2156 4132 2164
rect 4204 2156 4212 2164
rect 4108 2056 4116 2064
rect 4092 1956 4100 1964
rect 4204 2136 4212 2144
rect 4268 2136 4276 2144
rect 4316 2376 4324 2384
rect 4348 2336 4356 2344
rect 4316 2296 4324 2304
rect 4508 2676 4516 2684
rect 4508 2616 4516 2624
rect 4428 2596 4436 2604
rect 4476 2596 4484 2604
rect 4492 2596 4500 2604
rect 4476 2556 4484 2564
rect 4460 2516 4468 2524
rect 4444 2436 4452 2444
rect 4396 2396 4404 2404
rect 4428 2396 4436 2404
rect 4380 2336 4388 2344
rect 4348 2276 4356 2284
rect 4380 2276 4388 2284
rect 4252 2096 4260 2104
rect 4284 2096 4292 2104
rect 4316 2076 4324 2084
rect 4332 2076 4340 2084
rect 4156 2056 4164 2064
rect 4236 2056 4244 2064
rect 4268 2036 4276 2044
rect 4156 1996 4164 2004
rect 4108 1896 4116 1904
rect 4140 1896 4148 1904
rect 4172 1896 4180 1904
rect 4188 1896 4196 1904
rect 4236 1916 4244 1924
rect 4300 1956 4308 1964
rect 4204 1876 4212 1884
rect 4124 1856 4132 1864
rect 4092 1816 4100 1824
rect 4140 1816 4148 1824
rect 4108 1676 4116 1684
rect 4124 1676 4132 1684
rect 4268 1896 4276 1904
rect 4236 1796 4244 1804
rect 4220 1776 4228 1784
rect 4284 1796 4292 1804
rect 4188 1696 4196 1704
rect 4220 1676 4228 1684
rect 4140 1616 4148 1624
rect 4204 1576 4212 1584
rect 4124 1496 4132 1504
rect 3852 1476 3860 1484
rect 3932 1476 3940 1484
rect 3804 1436 3812 1444
rect 3900 1396 3908 1404
rect 3916 1396 3924 1404
rect 3932 1396 3940 1404
rect 3756 1376 3764 1384
rect 3676 1356 3684 1364
rect 3692 1316 3700 1324
rect 3676 1236 3684 1244
rect 3724 1216 3732 1224
rect 3804 1316 3812 1324
rect 3820 1236 3828 1244
rect 3724 1136 3732 1144
rect 3788 1136 3796 1144
rect 3836 1156 3844 1164
rect 3884 1156 3892 1164
rect 3756 1102 3764 1104
rect 3756 1096 3764 1102
rect 3852 1096 3860 1104
rect 3596 1036 3604 1044
rect 3628 1036 3636 1044
rect 3660 1036 3668 1044
rect 3612 996 3620 1004
rect 3644 996 3652 1004
rect 3484 956 3492 964
rect 3500 956 3508 964
rect 3564 956 3572 964
rect 3596 956 3604 964
rect 3532 916 3540 924
rect 3548 916 3556 924
rect 3468 896 3476 904
rect 3500 896 3508 904
rect 3516 896 3524 904
rect 3436 876 3444 884
rect 3420 756 3428 764
rect 3548 856 3556 864
rect 3692 976 3700 984
rect 3676 876 3684 884
rect 3644 856 3652 864
rect 3516 836 3524 844
rect 3564 836 3572 844
rect 3580 836 3588 844
rect 3372 716 3380 724
rect 3404 716 3412 724
rect 3324 636 3332 644
rect 3484 736 3492 744
rect 3500 736 3508 744
rect 3596 776 3604 784
rect 3660 776 3668 784
rect 3580 756 3588 764
rect 3436 676 3444 684
rect 3468 676 3476 684
rect 3372 596 3380 604
rect 3388 596 3396 604
rect 3452 616 3460 624
rect 3484 616 3492 624
rect 3516 716 3524 724
rect 3612 756 3620 764
rect 3612 716 3620 724
rect 3516 676 3524 684
rect 3644 696 3652 704
rect 3676 716 3684 724
rect 3612 656 3620 664
rect 3548 636 3556 644
rect 3580 636 3588 644
rect 3372 556 3380 564
rect 3196 456 3204 464
rect 3228 456 3236 464
rect 3148 396 3156 404
rect 3180 356 3188 364
rect 3132 316 3140 324
rect 3068 276 3076 284
rect 3084 276 3092 284
rect 3196 336 3204 344
rect 3196 316 3204 324
rect 2316 176 2324 184
rect 2348 176 2356 184
rect 2412 176 2420 184
rect 2428 176 2436 184
rect 2300 156 2308 164
rect 2332 156 2340 164
rect 2124 116 2132 124
rect 2204 116 2212 124
rect 2220 116 2228 124
rect 2236 116 2244 124
rect 2140 96 2148 104
rect 2172 96 2180 104
rect 2140 56 2148 64
rect 2156 56 2164 64
rect 2188 56 2196 64
rect 2204 56 2212 64
rect 140 16 148 24
rect 1548 16 1556 24
rect 1644 16 1652 24
rect 1577 6 1585 14
rect 1587 6 1595 14
rect 1597 6 1605 14
rect 1607 6 1615 14
rect 2140 16 2148 24
rect 2268 96 2276 104
rect 2284 96 2292 104
rect 2428 156 2436 164
rect 2460 156 2468 164
rect 2540 176 2548 184
rect 2444 136 2452 144
rect 2460 136 2468 144
rect 2492 136 2500 144
rect 2540 136 2548 144
rect 2476 116 2484 124
rect 2492 116 2500 124
rect 2364 96 2372 104
rect 2556 116 2564 124
rect 2620 116 2628 124
rect 2684 216 2692 224
rect 2764 196 2772 204
rect 2780 196 2788 204
rect 2812 216 2820 224
rect 2828 216 2836 224
rect 2812 196 2820 204
rect 2940 236 2948 244
rect 2956 236 2964 244
rect 2892 196 2900 204
rect 2396 96 2404 104
rect 2588 96 2596 104
rect 2508 76 2516 84
rect 2540 76 2548 84
rect 2364 56 2372 64
rect 2380 56 2388 64
rect 2380 36 2388 44
rect 2396 36 2404 44
rect 2556 36 2564 44
rect 2572 36 2580 44
rect 2620 36 2628 44
rect 3004 196 3012 204
rect 2972 156 2980 164
rect 2716 96 2724 104
rect 2732 96 2740 104
rect 2748 96 2756 104
rect 2812 96 2820 104
rect 2828 96 2836 104
rect 2732 76 2740 84
rect 2748 76 2756 84
rect 2796 76 2804 84
rect 2844 76 2852 84
rect 2668 36 2676 44
rect 2684 36 2692 44
rect 2764 56 2772 64
rect 2908 116 2916 124
rect 3052 256 3060 264
rect 3196 216 3204 224
rect 3113 206 3121 214
rect 3123 206 3131 214
rect 3133 206 3141 214
rect 3143 206 3151 214
rect 3084 196 3092 204
rect 2924 56 2932 64
rect 3324 536 3332 544
rect 3340 536 3348 544
rect 3324 516 3332 524
rect 3260 456 3268 464
rect 3228 336 3236 344
rect 3244 336 3252 344
rect 3356 516 3364 524
rect 3516 596 3524 604
rect 3420 536 3428 544
rect 3564 556 3572 564
rect 3580 556 3588 564
rect 3436 516 3444 524
rect 3500 536 3508 544
rect 3596 536 3604 544
rect 3516 516 3524 524
rect 3644 596 3652 604
rect 3660 576 3668 584
rect 3628 556 3636 564
rect 3676 556 3684 564
rect 3452 476 3460 484
rect 3324 376 3332 384
rect 3340 376 3348 384
rect 3292 336 3300 344
rect 3228 276 3236 284
rect 3276 276 3284 284
rect 3228 196 3236 204
rect 3244 176 3252 184
rect 3260 176 3268 184
rect 2860 36 2868 44
rect 2988 36 2996 44
rect 3036 36 3044 44
rect 3180 36 3188 44
rect 2716 16 2724 24
rect 2828 16 2836 24
rect 3228 96 3236 104
rect 3212 16 3220 24
rect 3324 336 3332 344
rect 3484 376 3492 384
rect 3420 336 3428 344
rect 3612 376 3620 384
rect 3532 336 3540 344
rect 3548 336 3556 344
rect 3580 336 3588 344
rect 3612 336 3620 344
rect 3340 276 3348 284
rect 3372 276 3380 284
rect 3340 236 3348 244
rect 3324 216 3332 224
rect 3308 176 3316 184
rect 3308 156 3316 164
rect 3324 156 3332 164
rect 3340 156 3348 164
rect 3308 136 3316 144
rect 3324 96 3332 104
rect 3420 216 3428 224
rect 3452 216 3460 224
rect 3484 276 3492 284
rect 3484 256 3492 264
rect 3468 156 3476 164
rect 3484 156 3492 164
rect 3468 136 3476 144
rect 3372 96 3380 104
rect 3452 36 3460 44
rect 3468 36 3476 44
rect 3516 316 3524 324
rect 3708 956 3716 964
rect 3804 1016 3812 1024
rect 4044 1416 4052 1424
rect 4108 1396 4116 1404
rect 4092 1356 4100 1364
rect 4012 1336 4020 1344
rect 4092 1336 4100 1344
rect 3980 1316 3988 1324
rect 4060 1316 4068 1324
rect 4012 1296 4020 1304
rect 3964 1236 3972 1244
rect 4028 1236 4036 1244
rect 3916 1196 3924 1204
rect 4092 1196 4100 1204
rect 4156 1416 4164 1424
rect 4188 1436 4196 1444
rect 4140 1396 4148 1404
rect 4172 1396 4180 1404
rect 4220 1376 4228 1384
rect 4172 1356 4180 1364
rect 4220 1316 4228 1324
rect 4044 1136 4052 1144
rect 3916 1116 3924 1124
rect 3900 1096 3908 1104
rect 3884 1056 3892 1064
rect 3996 1036 4004 1044
rect 3916 996 3924 1004
rect 3980 976 3988 984
rect 3740 936 3748 944
rect 3836 936 3844 944
rect 3708 896 3716 904
rect 3820 896 3828 904
rect 3740 796 3748 804
rect 3724 696 3732 704
rect 3820 756 3828 764
rect 3820 696 3828 704
rect 3788 676 3796 684
rect 3804 676 3812 684
rect 3692 496 3700 504
rect 3708 496 3716 504
rect 3708 416 3716 424
rect 3676 336 3684 344
rect 3740 656 3748 664
rect 3740 596 3748 604
rect 3772 596 3780 604
rect 3788 596 3796 604
rect 3756 576 3764 584
rect 3740 556 3748 564
rect 3756 556 3764 564
rect 3788 556 3796 564
rect 3852 856 3860 864
rect 3852 816 3860 824
rect 4172 1116 4180 1124
rect 4124 976 4132 984
rect 4156 976 4164 984
rect 4108 956 4116 964
rect 3900 936 3908 944
rect 3980 936 3988 944
rect 3916 816 3924 824
rect 3884 796 3892 804
rect 3868 776 3876 784
rect 3916 716 3924 724
rect 3900 696 3908 704
rect 3852 656 3860 664
rect 3836 636 3844 644
rect 3836 576 3844 584
rect 3820 556 3828 564
rect 3740 536 3748 544
rect 3804 536 3812 544
rect 3772 516 3780 524
rect 3884 596 3892 604
rect 3868 576 3876 584
rect 3868 496 3876 504
rect 3788 436 3796 444
rect 3820 396 3828 404
rect 3788 356 3796 364
rect 3804 356 3812 364
rect 3644 316 3652 324
rect 3708 316 3716 324
rect 3724 316 3732 324
rect 3596 276 3604 284
rect 3516 256 3524 264
rect 3564 256 3572 264
rect 3692 276 3700 284
rect 3708 196 3716 204
rect 3660 176 3668 184
rect 3708 156 3716 164
rect 3532 136 3540 144
rect 3516 116 3524 124
rect 3740 216 3748 224
rect 3996 816 4004 824
rect 4028 816 4036 824
rect 4156 876 4164 884
rect 4140 836 4148 844
rect 4108 756 4116 764
rect 4188 1036 4196 1044
rect 4204 1036 4212 1044
rect 4188 956 4196 964
rect 4252 1656 4260 1664
rect 4252 1616 4260 1624
rect 4252 1536 4260 1544
rect 4268 1536 4276 1544
rect 4364 2256 4372 2264
rect 4380 2176 4388 2184
rect 4364 2116 4372 2124
rect 4412 2336 4420 2344
rect 4428 2256 4436 2264
rect 4476 2476 4484 2484
rect 4508 2556 4516 2564
rect 4588 2676 4596 2684
rect 4540 2496 4548 2504
rect 4476 2396 4484 2404
rect 4665 2806 4673 2814
rect 4675 2806 4683 2814
rect 4685 2806 4693 2814
rect 4695 2806 4703 2814
rect 4796 2716 4804 2724
rect 4780 2696 4788 2704
rect 4844 2696 4852 2704
rect 5020 2696 5028 2704
rect 4860 2676 4868 2684
rect 4892 2676 4900 2684
rect 4908 2676 4916 2684
rect 4652 2656 4660 2664
rect 4764 2656 4772 2664
rect 4764 2596 4772 2604
rect 4652 2576 4660 2584
rect 4716 2576 4724 2584
rect 4652 2556 4660 2564
rect 4876 2656 4884 2664
rect 4972 2656 4980 2664
rect 4988 2576 4996 2584
rect 5020 2576 5028 2584
rect 4732 2536 4740 2544
rect 4860 2536 4868 2544
rect 4924 2536 4932 2544
rect 4572 2436 4580 2444
rect 4620 2436 4628 2444
rect 4524 2416 4532 2424
rect 4476 2336 4484 2344
rect 4524 2336 4532 2344
rect 4460 2276 4468 2284
rect 4444 2236 4452 2244
rect 4476 2236 4484 2244
rect 4476 2196 4484 2204
rect 4428 2176 4436 2184
rect 4508 2276 4516 2284
rect 4556 2236 4564 2244
rect 4572 2236 4580 2244
rect 4556 2196 4564 2204
rect 4492 2156 4500 2164
rect 4460 2136 4468 2144
rect 4476 2136 4484 2144
rect 4444 2116 4452 2124
rect 4556 2116 4564 2124
rect 4380 2096 4388 2104
rect 4396 2096 4404 2104
rect 4412 2056 4420 2064
rect 4428 1976 4436 1984
rect 4348 1956 4356 1964
rect 4332 1916 4340 1924
rect 4380 1896 4388 1904
rect 4332 1876 4340 1884
rect 4316 1796 4324 1804
rect 4460 1896 4468 1904
rect 4444 1876 4452 1884
rect 4380 1856 4388 1864
rect 4428 1856 4436 1864
rect 4316 1736 4324 1744
rect 4300 1656 4308 1664
rect 4316 1556 4324 1564
rect 4284 1476 4292 1484
rect 4252 1396 4260 1404
rect 4364 1756 4372 1764
rect 4412 1756 4420 1764
rect 4428 1736 4436 1744
rect 4380 1656 4388 1664
rect 4364 1576 4372 1584
rect 4364 1536 4372 1544
rect 4396 1516 4404 1524
rect 4348 1476 4356 1484
rect 4396 1456 4404 1464
rect 4508 2056 4516 2064
rect 4508 1956 4516 1964
rect 4588 2196 4596 2204
rect 4604 2196 4612 2204
rect 4588 2116 4596 2124
rect 4892 2496 4900 2504
rect 4748 2436 4756 2444
rect 4956 2496 4964 2504
rect 4665 2406 4673 2414
rect 4675 2406 4683 2414
rect 4685 2406 4693 2414
rect 4695 2406 4703 2414
rect 4668 2376 4676 2384
rect 4764 2376 4772 2384
rect 4748 2316 4756 2324
rect 4636 2276 4644 2284
rect 4652 2276 4660 2284
rect 4716 2276 4724 2284
rect 4636 2236 4644 2244
rect 4652 2236 4660 2244
rect 4620 2176 4628 2184
rect 4636 2176 4644 2184
rect 4716 2136 4724 2144
rect 4620 2116 4628 2124
rect 4700 2116 4708 2124
rect 4732 2116 4740 2124
rect 4604 2056 4612 2064
rect 4604 1936 4612 1944
rect 4572 1916 4580 1924
rect 4604 1916 4612 1924
rect 4540 1896 4548 1904
rect 4604 1896 4612 1904
rect 4556 1836 4564 1844
rect 4572 1816 4580 1824
rect 4524 1796 4532 1804
rect 4588 1796 4596 1804
rect 4444 1696 4452 1704
rect 4476 1696 4484 1704
rect 4572 1616 4580 1624
rect 4588 1616 4596 1624
rect 4460 1596 4468 1604
rect 4492 1596 4500 1604
rect 4428 1536 4436 1544
rect 4460 1456 4468 1464
rect 4412 1436 4420 1444
rect 4316 1376 4324 1384
rect 4396 1356 4404 1364
rect 4348 1336 4356 1344
rect 4268 1316 4276 1324
rect 4316 1296 4324 1304
rect 4316 1276 4324 1284
rect 4252 1236 4260 1244
rect 4300 1236 4308 1244
rect 4284 1156 4292 1164
rect 4396 1296 4404 1304
rect 4476 1296 4484 1304
rect 4348 1236 4356 1244
rect 4412 1236 4420 1244
rect 4380 1216 4388 1224
rect 4332 1176 4340 1184
rect 4332 1116 4340 1124
rect 4300 1096 4308 1104
rect 4412 1156 4420 1164
rect 4364 1096 4372 1104
rect 4380 1096 4388 1104
rect 4572 1576 4580 1584
rect 4508 1336 4516 1344
rect 4588 1476 4596 1484
rect 4556 1396 4564 1404
rect 4572 1376 4580 1384
rect 4492 1236 4500 1244
rect 4508 1236 4516 1244
rect 4460 1216 4468 1224
rect 4428 1076 4436 1084
rect 4332 1056 4340 1064
rect 4380 1056 4388 1064
rect 4268 976 4276 984
rect 4316 976 4324 984
rect 4220 916 4228 924
rect 4188 896 4196 904
rect 4220 896 4228 904
rect 4188 876 4196 884
rect 4060 716 4068 724
rect 4092 716 4100 724
rect 4140 716 4148 724
rect 4028 696 4036 704
rect 4044 696 4052 704
rect 3916 556 3924 564
rect 4108 656 4116 664
rect 4028 636 4036 644
rect 4092 636 4100 644
rect 3996 616 4004 624
rect 4012 616 4020 624
rect 3996 596 4004 604
rect 3980 576 3988 584
rect 4012 556 4020 564
rect 4028 536 4036 544
rect 4060 536 4068 544
rect 3932 496 3940 504
rect 3932 436 3940 444
rect 3900 416 3908 424
rect 3900 396 3908 404
rect 3884 356 3892 364
rect 3868 316 3876 324
rect 3916 376 3924 384
rect 3932 376 3940 384
rect 3916 276 3924 284
rect 3788 256 3796 264
rect 3804 256 3812 264
rect 3836 256 3844 264
rect 3756 196 3764 204
rect 3772 196 3780 204
rect 3804 156 3812 164
rect 3820 156 3828 164
rect 3580 136 3588 144
rect 3676 136 3684 144
rect 3724 136 3732 144
rect 3756 140 3764 144
rect 3756 136 3764 140
rect 3852 136 3860 144
rect 3676 116 3684 124
rect 3548 96 3556 104
rect 3644 96 3652 104
rect 3900 256 3908 264
rect 3964 496 3972 504
rect 3964 456 3972 464
rect 4044 436 4052 444
rect 4060 436 4068 444
rect 4060 376 4068 384
rect 4028 356 4036 364
rect 4092 356 4100 364
rect 3948 236 3956 244
rect 3964 216 3972 224
rect 3980 216 3988 224
rect 3916 156 3924 164
rect 4236 876 4244 884
rect 4204 736 4212 744
rect 4156 676 4164 684
rect 4204 716 4212 724
rect 4220 696 4228 704
rect 4204 676 4212 684
rect 4156 636 4164 644
rect 4140 596 4148 604
rect 4156 576 4164 584
rect 4364 1036 4372 1044
rect 4476 1036 4484 1044
rect 4540 1296 4548 1304
rect 4508 1176 4516 1184
rect 4524 1176 4532 1184
rect 4524 1136 4532 1144
rect 4556 1116 4564 1124
rect 4636 2056 4644 2064
rect 4636 2016 4644 2024
rect 4665 2006 4673 2014
rect 4675 2006 4683 2014
rect 4685 2006 4693 2014
rect 4695 2006 4703 2014
rect 4748 2076 4756 2084
rect 4892 2276 4900 2284
rect 4812 2256 4820 2264
rect 4860 2256 4868 2264
rect 4796 2236 4804 2244
rect 4828 2236 4836 2244
rect 4860 2236 4868 2244
rect 4780 2196 4788 2204
rect 4812 2176 4820 2184
rect 4764 2036 4772 2044
rect 4796 2036 4804 2044
rect 4828 2116 4836 2124
rect 4860 2116 4868 2124
rect 4876 2056 4884 2064
rect 4812 2016 4820 2024
rect 4652 1976 4660 1984
rect 4700 1976 4708 1984
rect 4732 1976 4740 1984
rect 4636 1936 4644 1944
rect 4652 1896 4660 1904
rect 4652 1796 4660 1804
rect 4988 2316 4996 2324
rect 5068 2916 5076 2924
rect 5500 3296 5508 3304
rect 5436 3276 5444 3284
rect 5468 3276 5476 3284
rect 5724 3476 5732 3484
rect 5724 3456 5732 3464
rect 5740 3436 5748 3444
rect 5820 3776 5828 3784
rect 5820 3676 5828 3684
rect 5836 3636 5844 3644
rect 5852 3616 5860 3624
rect 5852 3576 5860 3584
rect 5804 3536 5812 3544
rect 5772 3396 5780 3404
rect 5548 3356 5556 3364
rect 5596 3356 5604 3364
rect 5628 3356 5636 3364
rect 5644 3356 5652 3364
rect 5708 3356 5716 3364
rect 5740 3356 5748 3364
rect 5532 3316 5540 3324
rect 5596 3316 5604 3324
rect 5612 3316 5620 3324
rect 5580 3296 5588 3304
rect 5740 3336 5748 3344
rect 5660 3296 5668 3304
rect 5404 3196 5412 3204
rect 5836 3516 5844 3524
rect 5916 3856 5924 3864
rect 5900 3836 5908 3844
rect 5932 3756 5940 3764
rect 5884 3716 5892 3724
rect 5900 3716 5908 3724
rect 5884 3696 5892 3704
rect 5900 3656 5908 3664
rect 5932 3716 5940 3724
rect 6220 4316 6228 4324
rect 6172 4276 6180 4284
rect 6220 4276 6228 4284
rect 6188 4216 6196 4224
rect 6220 4216 6228 4224
rect 6156 4176 6164 4184
rect 6060 4076 6068 4084
rect 6092 4076 6100 4084
rect 6124 4076 6132 4084
rect 6060 4056 6068 4064
rect 5996 3976 6004 3984
rect 6028 3976 6036 3984
rect 6012 3956 6020 3964
rect 5996 3936 6004 3944
rect 5980 3916 5988 3924
rect 5964 3856 5972 3864
rect 5964 3736 5972 3744
rect 5916 3636 5924 3644
rect 5932 3616 5940 3624
rect 5868 3536 5876 3544
rect 5868 3516 5876 3524
rect 5900 3536 5908 3544
rect 5996 3876 6004 3884
rect 6140 4016 6148 4024
rect 6188 4156 6196 4164
rect 6268 4136 6276 4144
rect 6172 4116 6180 4124
rect 6220 4116 6228 4124
rect 6188 4096 6196 4104
rect 6220 4096 6228 4104
rect 6284 4096 6292 4104
rect 6220 4036 6228 4044
rect 6156 3996 6164 4004
rect 6076 3956 6084 3964
rect 6124 3916 6132 3924
rect 6108 3896 6116 3904
rect 6188 3896 6196 3904
rect 6028 3876 6036 3884
rect 6060 3876 6068 3884
rect 6220 3916 6228 3924
rect 6124 3876 6132 3884
rect 6012 3816 6020 3824
rect 5996 3796 6004 3804
rect 6044 3816 6052 3824
rect 6044 3776 6052 3784
rect 6188 3876 6196 3884
rect 6140 3856 6148 3864
rect 6156 3856 6164 3864
rect 6156 3836 6164 3844
rect 6172 3816 6180 3824
rect 6156 3796 6164 3804
rect 6092 3776 6100 3784
rect 6204 3856 6212 3864
rect 6028 3736 6036 3744
rect 5964 3616 5972 3624
rect 5980 3616 5988 3624
rect 5948 3576 5956 3584
rect 5980 3576 5988 3584
rect 5948 3536 5956 3544
rect 5852 3476 5860 3484
rect 5884 3476 5892 3484
rect 5932 3476 5940 3484
rect 5916 3416 5924 3424
rect 6044 3716 6052 3724
rect 6012 3636 6020 3644
rect 6028 3616 6036 3624
rect 6140 3716 6148 3724
rect 6156 3716 6164 3724
rect 6284 3936 6292 3944
rect 6220 3796 6228 3804
rect 6284 3836 6292 3844
rect 6252 3736 6260 3744
rect 6284 3736 6292 3744
rect 6124 3696 6132 3704
rect 6172 3696 6180 3704
rect 6188 3696 6196 3704
rect 6204 3696 6212 3704
rect 6236 3696 6244 3704
rect 6252 3696 6260 3704
rect 6108 3676 6116 3684
rect 5996 3516 6004 3524
rect 5964 3456 5972 3464
rect 5980 3436 5988 3444
rect 5948 3396 5956 3404
rect 5820 3376 5828 3384
rect 5820 3336 5828 3344
rect 5836 3336 5844 3344
rect 5804 3296 5812 3304
rect 5884 3336 5892 3344
rect 5900 3336 5908 3344
rect 5964 3336 5972 3344
rect 5900 3296 5908 3304
rect 5932 3296 5940 3304
rect 5996 3396 6004 3404
rect 6012 3376 6020 3384
rect 6092 3596 6100 3604
rect 6076 3556 6084 3564
rect 6044 3516 6052 3524
rect 6076 3476 6084 3484
rect 6076 3436 6084 3444
rect 6044 3416 6052 3424
rect 6028 3336 6036 3344
rect 6012 3316 6020 3324
rect 6028 3316 6036 3324
rect 5980 3296 5988 3304
rect 5948 3276 5956 3284
rect 5868 3256 5876 3264
rect 5164 3156 5172 3164
rect 5324 3156 5332 3164
rect 5756 3156 5764 3164
rect 5180 3116 5188 3124
rect 5276 3116 5284 3124
rect 5308 3116 5316 3124
rect 5212 3102 5220 3104
rect 5212 3096 5220 3102
rect 5276 3096 5284 3104
rect 5196 3056 5204 3064
rect 5292 3016 5300 3024
rect 5228 2996 5236 3004
rect 5260 2996 5268 3004
rect 5212 2956 5220 2964
rect 5148 2936 5156 2944
rect 5116 2896 5124 2904
rect 5196 2896 5204 2904
rect 5212 2896 5220 2904
rect 5116 2876 5124 2884
rect 5148 2716 5156 2724
rect 5068 2656 5076 2664
rect 5068 2396 5076 2404
rect 5068 2356 5076 2364
rect 5004 2236 5012 2244
rect 5036 2236 5044 2244
rect 5020 2196 5028 2204
rect 5004 2136 5012 2144
rect 5052 2136 5060 2144
rect 4732 1936 4740 1944
rect 4844 1936 4852 1944
rect 4876 1936 4884 1944
rect 4748 1896 4756 1904
rect 4764 1896 4772 1904
rect 4828 1896 4836 1904
rect 4860 1896 4868 1904
rect 4988 1976 4996 1984
rect 4924 1916 4932 1924
rect 4940 1916 4948 1924
rect 4860 1856 4868 1864
rect 4764 1836 4772 1844
rect 4716 1796 4724 1804
rect 4700 1776 4708 1784
rect 4684 1736 4692 1744
rect 4812 1816 4820 1824
rect 4892 1816 4900 1824
rect 5036 2096 5044 2104
rect 5036 2056 5044 2064
rect 5020 2016 5028 2024
rect 5100 2496 5108 2504
rect 5500 3136 5508 3144
rect 5596 3136 5604 3144
rect 5628 3136 5636 3144
rect 5420 3116 5428 3124
rect 5532 3116 5540 3124
rect 5596 3116 5604 3124
rect 5420 3096 5428 3104
rect 5452 3096 5460 3104
rect 5548 3096 5556 3104
rect 5324 3076 5332 3084
rect 5420 3076 5428 3084
rect 5452 3076 5460 3084
rect 5468 3076 5476 3084
rect 5516 3076 5524 3084
rect 5340 3056 5348 3064
rect 5404 3056 5412 3064
rect 5436 3056 5444 3064
rect 5388 3016 5396 3024
rect 5340 2956 5348 2964
rect 5372 2956 5380 2964
rect 5708 3096 5716 3104
rect 5804 3116 5812 3124
rect 5772 3076 5780 3084
rect 5836 3096 5844 3104
rect 5532 3036 5540 3044
rect 5676 3056 5684 3064
rect 5436 2956 5444 2964
rect 5516 2956 5524 2964
rect 5420 2936 5428 2944
rect 5276 2916 5284 2924
rect 5468 2876 5476 2884
rect 5548 2956 5556 2964
rect 5564 2956 5572 2964
rect 5516 2876 5524 2884
rect 5276 2856 5284 2864
rect 5324 2856 5332 2864
rect 5500 2856 5508 2864
rect 5500 2836 5508 2844
rect 5276 2776 5284 2784
rect 5468 2776 5476 2784
rect 5500 2736 5508 2744
rect 5516 2736 5524 2744
rect 5340 2716 5348 2724
rect 5244 2696 5252 2704
rect 5228 2676 5236 2684
rect 5308 2656 5316 2664
rect 5484 2656 5492 2664
rect 5292 2616 5300 2624
rect 5340 2616 5348 2624
rect 5500 2616 5508 2624
rect 5388 2596 5396 2604
rect 5484 2576 5492 2584
rect 5132 2536 5140 2544
rect 5324 2536 5332 2544
rect 5212 2496 5220 2504
rect 5260 2416 5268 2424
rect 5228 2396 5236 2404
rect 5244 2336 5252 2344
rect 5100 2296 5108 2304
rect 5084 2156 5092 2164
rect 5116 2136 5124 2144
rect 5100 2056 5108 2064
rect 5052 1936 5060 1944
rect 5084 1936 5092 1944
rect 5068 1896 5076 1904
rect 5436 2536 5444 2544
rect 5452 2536 5460 2544
rect 5644 2956 5652 2964
rect 5676 2996 5684 3004
rect 5724 3036 5732 3044
rect 5692 2976 5700 2984
rect 5836 3036 5844 3044
rect 5788 3016 5796 3024
rect 5804 2976 5812 2984
rect 5676 2956 5684 2964
rect 5740 2956 5748 2964
rect 5628 2916 5636 2924
rect 5580 2856 5588 2864
rect 5692 2936 5700 2944
rect 5740 2936 5748 2944
rect 5692 2896 5700 2904
rect 5724 2856 5732 2864
rect 5708 2836 5716 2844
rect 5676 2816 5684 2824
rect 5596 2796 5604 2804
rect 5628 2796 5636 2804
rect 5580 2736 5588 2744
rect 5564 2716 5572 2724
rect 5628 2716 5636 2724
rect 5788 2896 5796 2904
rect 5820 2876 5828 2884
rect 5724 2756 5732 2764
rect 5740 2756 5748 2764
rect 5804 2756 5812 2764
rect 5548 2636 5556 2644
rect 5772 2736 5780 2744
rect 5756 2696 5764 2704
rect 5804 2696 5812 2704
rect 5772 2676 5780 2684
rect 5804 2656 5812 2664
rect 5740 2616 5748 2624
rect 5788 2616 5796 2624
rect 5708 2596 5716 2604
rect 5756 2536 5764 2544
rect 5692 2516 5700 2524
rect 5804 2516 5812 2524
rect 5516 2496 5524 2504
rect 5628 2496 5636 2504
rect 5708 2496 5716 2504
rect 5788 2496 5796 2504
rect 5436 2476 5444 2484
rect 5756 2476 5764 2484
rect 5548 2436 5556 2444
rect 5612 2436 5620 2444
rect 5692 2436 5700 2444
rect 5724 2436 5732 2444
rect 5740 2436 5748 2444
rect 5612 2316 5620 2324
rect 5644 2316 5652 2324
rect 5276 2296 5284 2304
rect 5372 2296 5380 2304
rect 5580 2302 5588 2304
rect 5580 2296 5588 2302
rect 5644 2296 5652 2304
rect 5724 2416 5732 2424
rect 5420 2276 5428 2284
rect 5516 2276 5524 2284
rect 5676 2276 5684 2284
rect 5164 2216 5172 2224
rect 5180 2176 5188 2184
rect 5212 2136 5220 2144
rect 5148 2116 5156 2124
rect 5196 2036 5204 2044
rect 5164 1956 5172 1964
rect 5692 2256 5700 2264
rect 5676 2196 5684 2204
rect 5356 2136 5364 2144
rect 5500 2136 5508 2144
rect 5676 2136 5684 2144
rect 5260 2116 5268 2124
rect 5324 2118 5332 2124
rect 5324 2116 5332 2118
rect 5356 2116 5364 2124
rect 5420 2116 5428 2124
rect 5468 2116 5476 2124
rect 5324 2076 5332 2084
rect 5324 2056 5332 2064
rect 5196 1936 5204 1944
rect 5228 1936 5236 1944
rect 5244 1936 5252 1944
rect 5340 1936 5348 1944
rect 5388 2056 5396 2064
rect 5404 1936 5412 1944
rect 5564 1936 5572 1944
rect 5372 1896 5380 1904
rect 5436 1896 5444 1904
rect 5084 1876 5092 1884
rect 5148 1876 5156 1884
rect 5132 1856 5140 1864
rect 5116 1816 5124 1824
rect 4988 1776 4996 1784
rect 5052 1776 5060 1784
rect 4716 1696 4724 1704
rect 4796 1696 4804 1704
rect 4652 1656 4660 1664
rect 4812 1656 4820 1664
rect 4876 1656 4884 1664
rect 4860 1636 4868 1644
rect 4844 1616 4852 1624
rect 4665 1606 4673 1614
rect 4675 1606 4683 1614
rect 4685 1606 4693 1614
rect 4695 1606 4703 1614
rect 4636 1596 4644 1604
rect 4732 1596 4740 1604
rect 4668 1576 4676 1584
rect 4684 1576 4692 1584
rect 4860 1536 4868 1544
rect 4732 1516 4740 1524
rect 4764 1516 4772 1524
rect 4828 1516 4836 1524
rect 4636 1476 4644 1484
rect 4812 1476 4820 1484
rect 4828 1476 4836 1484
rect 4668 1456 4676 1464
rect 4620 1396 4628 1404
rect 4604 1116 4612 1124
rect 4620 1096 4628 1104
rect 4540 1016 4548 1024
rect 4492 976 4500 984
rect 4348 956 4356 964
rect 4508 916 4516 924
rect 4604 976 4612 984
rect 4652 1396 4660 1404
rect 4716 1436 4724 1444
rect 4668 1376 4676 1384
rect 4652 1336 4660 1344
rect 4780 1396 4788 1404
rect 4828 1396 4836 1404
rect 4876 1516 4884 1524
rect 4972 1736 4980 1744
rect 5036 1736 5044 1744
rect 5068 1736 5076 1744
rect 5084 1736 5092 1744
rect 4924 1676 4932 1684
rect 4908 1656 4916 1664
rect 5004 1636 5012 1644
rect 4956 1616 4964 1624
rect 4956 1516 4964 1524
rect 4860 1436 4868 1444
rect 4844 1376 4852 1384
rect 4860 1376 4868 1384
rect 4748 1336 4756 1344
rect 4716 1276 4724 1284
rect 4665 1206 4673 1214
rect 4675 1206 4683 1214
rect 4685 1206 4693 1214
rect 4695 1206 4703 1214
rect 4732 1176 4740 1184
rect 4668 1156 4676 1164
rect 4652 1116 4660 1124
rect 4652 1036 4660 1044
rect 4348 896 4356 904
rect 4396 896 4404 904
rect 4412 896 4420 904
rect 4476 896 4484 904
rect 4572 916 4580 924
rect 4636 916 4644 924
rect 4284 876 4292 884
rect 4348 876 4356 884
rect 4332 796 4340 804
rect 4300 716 4308 724
rect 4268 676 4276 684
rect 4364 816 4372 824
rect 4380 796 4388 804
rect 4348 716 4356 724
rect 4220 636 4228 644
rect 4268 616 4276 624
rect 4172 556 4180 564
rect 4204 556 4212 564
rect 4124 536 4132 544
rect 4204 536 4212 544
rect 4140 476 4148 484
rect 4156 356 4164 364
rect 4172 356 4180 364
rect 4060 282 4068 284
rect 4060 276 4068 282
rect 4092 296 4100 304
rect 4108 296 4116 304
rect 4252 496 4260 504
rect 4300 576 4308 584
rect 4284 556 4292 564
rect 4316 556 4324 564
rect 4268 476 4276 484
rect 4284 476 4292 484
rect 4220 396 4228 404
rect 4204 376 4212 384
rect 4236 376 4244 384
rect 4188 336 4196 344
rect 4028 216 4036 224
rect 4140 236 4148 244
rect 3884 116 3892 124
rect 3852 96 3860 104
rect 3868 96 3876 104
rect 3900 96 3908 104
rect 3948 96 3956 104
rect 3676 56 3684 64
rect 4140 176 4148 184
rect 4156 156 4164 164
rect 4188 156 4196 164
rect 4108 136 4116 144
rect 4124 136 4132 144
rect 3980 76 3988 84
rect 4044 96 4052 104
rect 4092 96 4100 104
rect 4188 96 4196 104
rect 4028 76 4036 84
rect 4124 76 4132 84
rect 4220 176 4228 184
rect 4268 356 4276 364
rect 4252 276 4260 284
rect 4364 676 4372 684
rect 4380 676 4388 684
rect 4348 516 4356 524
rect 4332 496 4340 504
rect 4316 416 4324 424
rect 4332 356 4340 364
rect 4428 876 4436 884
rect 4540 876 4548 884
rect 4412 816 4420 824
rect 4620 896 4628 904
rect 4636 896 4644 904
rect 4588 836 4596 844
rect 4508 816 4516 824
rect 4460 796 4468 804
rect 4492 796 4500 804
rect 4444 776 4452 784
rect 4428 716 4436 724
rect 4460 716 4468 724
rect 4492 716 4500 724
rect 4524 796 4532 804
rect 4572 816 4580 824
rect 4604 716 4612 724
rect 4620 716 4628 724
rect 4844 1316 4852 1324
rect 4764 1296 4772 1304
rect 4780 1216 4788 1224
rect 4732 1096 4740 1104
rect 4828 1176 4836 1184
rect 4796 1136 4804 1144
rect 4860 1296 4868 1304
rect 4908 1476 4916 1484
rect 4940 1476 4948 1484
rect 4892 1416 4900 1424
rect 5020 1536 5028 1544
rect 5020 1496 5028 1504
rect 5068 1636 5076 1644
rect 5308 1876 5316 1884
rect 5388 1876 5396 1884
rect 5260 1856 5268 1864
rect 5452 1856 5460 1864
rect 5500 1856 5508 1864
rect 5244 1816 5252 1824
rect 5436 1776 5444 1784
rect 5260 1736 5268 1744
rect 5484 1816 5492 1824
rect 5500 1816 5508 1824
rect 5468 1756 5476 1764
rect 5468 1736 5476 1744
rect 5532 1776 5540 1784
rect 5516 1756 5524 1764
rect 5532 1756 5540 1764
rect 5196 1696 5204 1704
rect 5148 1656 5156 1664
rect 5084 1616 5092 1624
rect 5068 1496 5076 1504
rect 5036 1476 5044 1484
rect 4988 1396 4996 1404
rect 4924 1376 4932 1384
rect 4956 1356 4964 1364
rect 5004 1356 5012 1364
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 4892 1296 4900 1304
rect 4924 1296 4932 1304
rect 4940 1296 4948 1304
rect 4972 1236 4980 1244
rect 4876 1136 4884 1144
rect 4908 1136 4916 1144
rect 4812 1096 4820 1104
rect 4796 1036 4804 1044
rect 4700 1016 4708 1024
rect 4780 1016 4788 1024
rect 4668 876 4676 884
rect 4732 916 4740 924
rect 4780 896 4788 904
rect 4764 876 4772 884
rect 4665 806 4673 814
rect 4675 806 4683 814
rect 4685 806 4693 814
rect 4695 806 4703 814
rect 4668 776 4676 784
rect 4556 676 4564 684
rect 4604 676 4612 684
rect 4412 656 4420 664
rect 4572 656 4580 664
rect 4412 596 4420 604
rect 4460 616 4468 624
rect 4524 636 4532 644
rect 4572 636 4580 644
rect 4588 636 4596 644
rect 4444 476 4452 484
rect 4396 416 4404 424
rect 4428 336 4436 344
rect 4300 276 4308 284
rect 4364 276 4372 284
rect 4268 156 4276 164
rect 4236 96 4244 104
rect 4284 136 4292 144
rect 4332 236 4340 244
rect 4428 256 4436 264
rect 4380 216 4388 224
rect 4380 176 4388 184
rect 4316 116 4324 124
rect 4364 156 4372 164
rect 4412 156 4420 164
rect 4492 576 4500 584
rect 4748 816 4756 824
rect 4732 736 4740 744
rect 4764 716 4772 724
rect 4764 676 4772 684
rect 4876 1076 4884 1084
rect 4844 1036 4852 1044
rect 4940 1136 4948 1144
rect 5020 1296 5028 1304
rect 5052 1416 5060 1424
rect 5100 1416 5108 1424
rect 5052 1376 5060 1384
rect 5052 1356 5060 1364
rect 5020 1256 5028 1264
rect 5036 1256 5044 1264
rect 5004 1136 5012 1144
rect 4988 1096 4996 1104
rect 5276 1696 5284 1704
rect 5292 1696 5300 1704
rect 5388 1696 5396 1704
rect 5532 1696 5540 1704
rect 5436 1676 5444 1684
rect 5276 1616 5284 1624
rect 5260 1556 5268 1564
rect 5212 1516 5220 1524
rect 5292 1516 5300 1524
rect 5308 1516 5316 1524
rect 5340 1516 5348 1524
rect 5244 1496 5252 1504
rect 5244 1456 5252 1464
rect 5292 1456 5300 1464
rect 5196 1356 5204 1364
rect 5132 1316 5140 1324
rect 5068 1256 5076 1264
rect 5132 1296 5140 1304
rect 5084 1236 5092 1244
rect 5068 1216 5076 1224
rect 4972 1076 4980 1084
rect 5004 1076 5012 1084
rect 4828 756 4836 764
rect 4828 716 4836 724
rect 4892 976 4900 984
rect 4908 976 4916 984
rect 4924 976 4932 984
rect 4892 916 4900 924
rect 4876 896 4884 904
rect 5052 1076 5060 1084
rect 5148 1216 5156 1224
rect 5180 1176 5188 1184
rect 5132 1156 5140 1164
rect 5100 1136 5108 1144
rect 5116 1116 5124 1124
rect 5180 1116 5188 1124
rect 5100 1076 5108 1084
rect 5116 1076 5124 1084
rect 5148 1076 5156 1084
rect 4892 876 4900 884
rect 4908 876 4916 884
rect 4988 1036 4996 1044
rect 5052 1036 5060 1044
rect 4972 1016 4980 1024
rect 5036 1016 5044 1024
rect 4988 976 4996 984
rect 5020 976 5028 984
rect 5020 916 5028 924
rect 4956 876 4964 884
rect 4908 776 4916 784
rect 4956 796 4964 804
rect 4940 756 4948 764
rect 4652 636 4660 644
rect 4540 516 4548 524
rect 4492 496 4500 504
rect 4508 436 4516 444
rect 4476 396 4484 404
rect 4492 396 4500 404
rect 4524 396 4532 404
rect 4460 356 4468 364
rect 4652 576 4660 584
rect 4604 536 4612 544
rect 4620 536 4628 544
rect 4588 456 4596 464
rect 4556 396 4564 404
rect 4556 356 4564 364
rect 4492 336 4500 344
rect 4540 336 4548 344
rect 4508 316 4516 324
rect 4476 296 4484 304
rect 4812 656 4820 664
rect 4764 636 4772 644
rect 4700 496 4708 504
rect 4700 456 4708 464
rect 4636 436 4644 444
rect 4684 436 4692 444
rect 4604 396 4612 404
rect 4604 376 4612 384
rect 4620 356 4628 364
rect 4604 336 4612 344
rect 4460 256 4468 264
rect 4492 256 4500 264
rect 4588 276 4596 284
rect 4460 236 4468 244
rect 4665 406 4673 414
rect 4675 406 4683 414
rect 4685 406 4693 414
rect 4695 406 4703 414
rect 4732 396 4740 404
rect 4748 376 4756 384
rect 4732 336 4740 344
rect 4796 576 4804 584
rect 4796 516 4804 524
rect 4812 516 4820 524
rect 5020 876 5028 884
rect 5004 756 5012 764
rect 4972 716 4980 724
rect 5020 716 5028 724
rect 5084 1016 5092 1024
rect 5052 916 5060 924
rect 5068 876 5076 884
rect 5068 836 5076 844
rect 5148 956 5156 964
rect 5100 916 5108 924
rect 5100 876 5108 884
rect 5116 876 5124 884
rect 5068 816 5076 824
rect 5084 816 5092 824
rect 5132 816 5140 824
rect 5148 816 5156 824
rect 5404 1476 5412 1484
rect 5420 1476 5428 1484
rect 5324 1456 5332 1464
rect 5420 1456 5428 1464
rect 5308 1416 5316 1424
rect 5340 1356 5348 1364
rect 5276 1336 5284 1344
rect 5308 1316 5316 1324
rect 5212 1276 5220 1284
rect 5292 1276 5300 1284
rect 5308 1276 5316 1284
rect 5212 1216 5220 1224
rect 5372 1316 5380 1324
rect 5404 1256 5412 1264
rect 5340 1236 5348 1244
rect 5308 1216 5316 1224
rect 5340 1156 5348 1164
rect 5292 1136 5300 1144
rect 5276 1116 5284 1124
rect 5372 1116 5380 1124
rect 5372 1096 5380 1104
rect 5308 1076 5316 1084
rect 5372 1076 5380 1084
rect 5452 1656 5460 1664
rect 5612 2016 5620 2024
rect 5596 1936 5604 1944
rect 5580 1916 5588 1924
rect 5660 1916 5668 1924
rect 5612 1816 5620 1824
rect 5676 1876 5684 1884
rect 5708 2196 5716 2204
rect 5708 1976 5716 1984
rect 5772 2376 5780 2384
rect 5740 2296 5748 2304
rect 5948 3236 5956 3244
rect 5948 3176 5956 3184
rect 5900 3156 5908 3164
rect 5916 3136 5924 3144
rect 5964 3156 5972 3164
rect 5884 3116 5892 3124
rect 5900 3116 5908 3124
rect 5916 3096 5924 3104
rect 5884 3076 5892 3084
rect 5932 3076 5940 3084
rect 5868 2996 5876 3004
rect 5996 3156 6004 3164
rect 5980 3136 5988 3144
rect 5980 3096 5988 3104
rect 6140 3556 6148 3564
rect 6156 3456 6164 3464
rect 6124 3436 6132 3444
rect 6092 3416 6100 3424
rect 6060 3396 6068 3404
rect 6172 3376 6180 3384
rect 6140 3356 6148 3364
rect 6060 3336 6068 3344
rect 6076 3296 6084 3304
rect 6028 3256 6036 3264
rect 6044 3256 6052 3264
rect 6044 3176 6052 3184
rect 6028 3156 6036 3164
rect 5980 3056 5988 3064
rect 5980 2956 5988 2964
rect 5964 2896 5972 2904
rect 5996 2896 6004 2904
rect 5884 2856 5892 2864
rect 5868 2816 5876 2824
rect 5852 2776 5860 2784
rect 5884 2756 5892 2764
rect 5900 2736 5908 2744
rect 5868 2716 5876 2724
rect 5932 2716 5940 2724
rect 5948 2716 5956 2724
rect 5868 2676 5876 2684
rect 5932 2636 5940 2644
rect 5852 2616 5860 2624
rect 5900 2616 5908 2624
rect 5836 2536 5844 2544
rect 6108 3276 6116 3284
rect 6140 3296 6148 3304
rect 6108 3256 6116 3264
rect 6092 3176 6100 3184
rect 6092 3156 6100 3164
rect 6060 3116 6068 3124
rect 6124 3116 6132 3124
rect 6044 3056 6052 3064
rect 6076 3056 6084 3064
rect 6044 3036 6052 3044
rect 6076 2956 6084 2964
rect 6028 2936 6036 2944
rect 6060 2936 6068 2944
rect 6076 2936 6084 2944
rect 6012 2876 6020 2884
rect 5996 2856 6004 2864
rect 6028 2856 6036 2864
rect 5980 2736 5988 2744
rect 5980 2656 5988 2664
rect 5964 2636 5972 2644
rect 6012 2796 6020 2804
rect 6012 2656 6020 2664
rect 6028 2656 6036 2664
rect 6044 2636 6052 2644
rect 5996 2616 6004 2624
rect 6012 2596 6020 2604
rect 5996 2556 6004 2564
rect 5964 2536 5972 2544
rect 5916 2496 5924 2504
rect 5964 2516 5972 2524
rect 6028 2516 6036 2524
rect 5932 2456 5940 2464
rect 5900 2416 5908 2424
rect 5804 2296 5812 2304
rect 5916 2276 5924 2284
rect 5948 2276 5956 2284
rect 5804 2236 5812 2244
rect 5948 2236 5956 2244
rect 5820 2196 5828 2204
rect 5868 2196 5876 2204
rect 5820 2156 5828 2164
rect 5852 2156 5860 2164
rect 5820 2116 5828 2124
rect 5852 2116 5860 2124
rect 5868 2116 5876 2124
rect 5772 2016 5780 2024
rect 5916 2096 5924 2104
rect 5836 2076 5844 2084
rect 5804 1976 5812 1984
rect 5740 1956 5748 1964
rect 5932 1956 5940 1964
rect 5820 1916 5828 1924
rect 5772 1876 5780 1884
rect 5612 1776 5620 1784
rect 5644 1776 5652 1784
rect 5580 1756 5588 1764
rect 5596 1756 5604 1764
rect 5628 1716 5636 1724
rect 5612 1696 5620 1704
rect 5596 1676 5604 1684
rect 5580 1656 5588 1664
rect 5612 1656 5620 1664
rect 5564 1636 5572 1644
rect 5596 1636 5604 1644
rect 5468 1576 5476 1584
rect 5500 1516 5508 1524
rect 5548 1516 5556 1524
rect 5452 1416 5460 1424
rect 5532 1496 5540 1504
rect 5548 1476 5556 1484
rect 5660 1696 5668 1704
rect 5724 1856 5732 1864
rect 5724 1836 5732 1844
rect 5900 1836 5908 1844
rect 5868 1796 5876 1804
rect 5788 1776 5796 1784
rect 5724 1756 5732 1764
rect 5868 1756 5876 1764
rect 5820 1736 5828 1744
rect 5692 1716 5700 1724
rect 5724 1716 5732 1724
rect 5836 1716 5844 1724
rect 5660 1576 5668 1584
rect 5676 1496 5684 1504
rect 5644 1436 5652 1444
rect 5628 1376 5636 1384
rect 5532 1336 5540 1344
rect 5532 1316 5540 1324
rect 5516 1196 5524 1204
rect 5484 1136 5492 1144
rect 5420 1076 5428 1084
rect 5244 1036 5252 1044
rect 5308 1036 5316 1044
rect 5324 1036 5332 1044
rect 5372 1036 5380 1044
rect 5404 1036 5412 1044
rect 5276 996 5284 1004
rect 5212 956 5220 964
rect 5356 956 5364 964
rect 5196 936 5204 944
rect 5324 936 5332 944
rect 5340 936 5348 944
rect 5212 916 5220 924
rect 5276 916 5284 924
rect 5308 916 5316 924
rect 5068 756 5076 764
rect 5100 756 5108 764
rect 5132 756 5140 764
rect 5164 756 5172 764
rect 4972 656 4980 664
rect 4924 636 4932 644
rect 4956 636 4964 644
rect 4876 616 4884 624
rect 4940 616 4948 624
rect 4908 576 4916 584
rect 4924 576 4932 584
rect 4988 596 4996 604
rect 4876 556 4884 564
rect 4924 516 4932 524
rect 4860 496 4868 504
rect 4796 396 4804 404
rect 4860 396 4868 404
rect 4476 156 4484 164
rect 4604 236 4612 244
rect 4636 236 4644 244
rect 4588 216 4596 224
rect 4556 176 4564 184
rect 4380 116 4388 124
rect 4444 116 4452 124
rect 4332 56 4340 64
rect 4204 36 4212 44
rect 4492 96 4500 104
rect 4492 76 4500 84
rect 4412 56 4420 64
rect 4604 196 4612 204
rect 4620 176 4628 184
rect 4588 116 4596 124
rect 4684 216 4692 224
rect 4668 196 4676 204
rect 4540 56 4548 64
rect 4668 36 4676 44
rect 3356 16 3364 24
rect 3500 16 3508 24
rect 4636 16 4644 24
rect 4665 6 4673 14
rect 4675 6 4683 14
rect 4685 6 4693 14
rect 4695 6 4703 14
rect 4764 276 4772 284
rect 4828 376 4836 384
rect 4844 356 4852 364
rect 4812 296 4820 304
rect 4828 296 4836 304
rect 4748 236 4756 244
rect 4764 216 4772 224
rect 4780 216 4788 224
rect 4812 196 4820 204
rect 4908 476 4916 484
rect 4892 416 4900 424
rect 4940 456 4948 464
rect 4876 296 4884 304
rect 4860 276 4868 284
rect 4876 216 4884 224
rect 4876 196 4884 204
rect 4780 116 4788 124
rect 4796 116 4804 124
rect 4828 116 4836 124
rect 4748 36 4756 44
rect 5052 636 5060 644
rect 5004 576 5012 584
rect 5036 596 5044 604
rect 4988 496 4996 504
rect 4956 396 4964 404
rect 4956 296 4964 304
rect 5148 716 5156 724
rect 5148 656 5156 664
rect 5116 596 5124 604
rect 5260 896 5268 904
rect 5292 896 5300 904
rect 5244 876 5252 884
rect 5244 696 5252 704
rect 5244 656 5252 664
rect 5228 616 5236 624
rect 5212 596 5220 604
rect 5196 576 5204 584
rect 5084 516 5092 524
rect 5020 456 5028 464
rect 5036 416 5044 424
rect 5116 516 5124 524
rect 5180 516 5188 524
rect 5132 456 5140 464
rect 5148 396 5156 404
rect 5100 376 5108 384
rect 5068 356 5076 364
rect 5084 356 5092 364
rect 5164 376 5172 384
rect 5052 336 5060 344
rect 5004 316 5012 324
rect 5068 316 5076 324
rect 5020 296 5028 304
rect 4956 256 4964 264
rect 5020 256 5028 264
rect 5116 316 5124 324
rect 5100 296 5108 304
rect 4988 236 4996 244
rect 4972 216 4980 224
rect 5036 216 5044 224
rect 5020 176 5028 184
rect 5084 176 5092 184
rect 5052 156 5060 164
rect 4924 116 4932 124
rect 4940 116 4948 124
rect 5116 256 5124 264
rect 5324 876 5332 884
rect 5436 1056 5444 1064
rect 5420 996 5428 1004
rect 5436 996 5444 1004
rect 5532 1096 5540 1104
rect 5580 1256 5588 1264
rect 5580 1236 5588 1244
rect 5596 1196 5604 1204
rect 5564 1156 5572 1164
rect 5532 1076 5540 1084
rect 5548 1076 5556 1084
rect 5484 1036 5492 1044
rect 5500 1036 5508 1044
rect 5516 1016 5524 1024
rect 5516 996 5524 1004
rect 5468 976 5476 984
rect 5388 956 5396 964
rect 5596 1136 5604 1144
rect 5676 1416 5684 1424
rect 5676 1336 5684 1344
rect 5708 1676 5716 1684
rect 5804 1656 5812 1664
rect 5836 1656 5844 1664
rect 5868 1636 5876 1644
rect 5884 1636 5892 1644
rect 5836 1596 5844 1604
rect 5804 1576 5812 1584
rect 5756 1556 5764 1564
rect 5820 1556 5828 1564
rect 5836 1556 5844 1564
rect 5756 1516 5764 1524
rect 5740 1496 5748 1504
rect 5804 1496 5812 1504
rect 5772 1476 5780 1484
rect 5724 1456 5732 1464
rect 5708 1336 5716 1344
rect 5724 1296 5732 1304
rect 5724 1276 5732 1284
rect 5692 1256 5700 1264
rect 5676 1176 5684 1184
rect 5676 1156 5684 1164
rect 5580 1096 5588 1104
rect 5628 1096 5636 1104
rect 5532 956 5540 964
rect 5420 936 5428 944
rect 5436 936 5444 944
rect 5500 936 5508 944
rect 5308 816 5316 824
rect 5276 776 5284 784
rect 5276 756 5284 764
rect 5372 776 5380 784
rect 5260 616 5268 624
rect 5340 656 5348 664
rect 5356 636 5364 644
rect 5452 916 5460 924
rect 5468 916 5476 924
rect 5500 916 5508 924
rect 5532 916 5540 924
rect 5436 896 5444 904
rect 5468 876 5476 884
rect 5484 876 5492 884
rect 5436 856 5444 864
rect 5452 856 5460 864
rect 5436 816 5444 824
rect 5420 656 5428 664
rect 5260 556 5268 564
rect 5244 516 5252 524
rect 5212 476 5220 484
rect 5228 476 5236 484
rect 5228 456 5236 464
rect 5196 376 5204 384
rect 5180 316 5188 324
rect 5212 316 5220 324
rect 5164 256 5172 264
rect 5340 596 5348 604
rect 5372 616 5380 624
rect 5420 576 5428 584
rect 5372 556 5380 564
rect 5420 536 5428 544
rect 5420 516 5428 524
rect 5388 496 5396 504
rect 5340 476 5348 484
rect 5276 456 5284 464
rect 5340 416 5348 424
rect 5260 356 5268 364
rect 5276 336 5284 344
rect 5196 236 5204 244
rect 5228 236 5236 244
rect 5244 236 5252 244
rect 5212 196 5220 204
rect 5148 176 5156 184
rect 5180 176 5188 184
rect 5148 156 5156 164
rect 5116 136 5124 144
rect 5132 136 5140 144
rect 5068 116 5076 124
rect 5084 116 5092 124
rect 4940 76 4948 84
rect 5180 116 5188 124
rect 5244 116 5252 124
rect 5276 236 5284 244
rect 5372 356 5380 364
rect 5372 316 5380 324
rect 5356 296 5364 304
rect 5340 216 5348 224
rect 5324 176 5332 184
rect 5308 136 5316 144
rect 5468 776 5476 784
rect 5468 756 5476 764
rect 5564 1016 5572 1024
rect 5628 1056 5636 1064
rect 5612 1036 5620 1044
rect 5628 1036 5636 1044
rect 5612 996 5620 1004
rect 5580 956 5588 964
rect 5612 956 5620 964
rect 5628 956 5636 964
rect 5596 936 5604 944
rect 5612 936 5620 944
rect 5564 916 5572 924
rect 5548 896 5556 904
rect 5548 876 5556 884
rect 5516 856 5524 864
rect 5500 696 5508 704
rect 5532 756 5540 764
rect 5564 856 5572 864
rect 5660 1096 5668 1104
rect 5660 956 5668 964
rect 5740 1136 5748 1144
rect 5692 1096 5700 1104
rect 5708 1096 5716 1104
rect 5708 1076 5716 1084
rect 5724 1076 5732 1084
rect 5724 1016 5732 1024
rect 5692 956 5700 964
rect 5708 956 5716 964
rect 5788 1456 5796 1464
rect 5804 1396 5812 1404
rect 5804 1316 5812 1324
rect 5772 1136 5780 1144
rect 5836 1476 5844 1484
rect 5852 1476 5860 1484
rect 5836 1376 5844 1384
rect 5820 1216 5828 1224
rect 5868 1196 5876 1204
rect 5836 1136 5844 1144
rect 5788 1096 5796 1104
rect 5772 1076 5780 1084
rect 5804 1076 5812 1084
rect 5820 1076 5828 1084
rect 5756 1056 5764 1064
rect 5772 1036 5780 1044
rect 5740 956 5748 964
rect 5644 916 5652 924
rect 5676 916 5684 924
rect 5612 856 5620 864
rect 5628 856 5636 864
rect 5660 856 5668 864
rect 5628 836 5636 844
rect 5596 776 5604 784
rect 5612 776 5620 784
rect 5644 816 5652 824
rect 5708 936 5716 944
rect 5724 936 5732 944
rect 5820 1036 5828 1044
rect 5676 836 5684 844
rect 5692 836 5700 844
rect 5452 656 5460 664
rect 5436 496 5444 504
rect 5420 476 5428 484
rect 5564 656 5572 664
rect 5468 616 5476 624
rect 5548 616 5556 624
rect 5724 916 5732 924
rect 5804 936 5812 944
rect 5804 916 5812 924
rect 5788 896 5796 904
rect 5740 876 5748 884
rect 5804 816 5812 824
rect 5724 796 5732 804
rect 5692 776 5700 784
rect 5708 776 5716 784
rect 5740 756 5748 764
rect 5804 756 5812 764
rect 5692 696 5700 704
rect 5596 636 5604 644
rect 5644 636 5652 644
rect 5676 636 5684 644
rect 5564 596 5572 604
rect 5484 536 5492 544
rect 5516 556 5524 564
rect 5468 496 5476 504
rect 5452 416 5460 424
rect 5500 496 5508 504
rect 5500 476 5508 484
rect 5500 416 5508 424
rect 5548 536 5556 544
rect 5580 536 5588 544
rect 5628 616 5636 624
rect 5676 596 5684 604
rect 5756 636 5764 644
rect 5868 1176 5876 1184
rect 6044 2496 6052 2504
rect 6044 2476 6052 2484
rect 6076 2716 6084 2724
rect 6076 2636 6084 2644
rect 6076 2556 6084 2564
rect 6156 3136 6164 3144
rect 6156 3116 6164 3124
rect 6156 3096 6164 3104
rect 6108 3056 6116 3064
rect 6140 3056 6148 3064
rect 6156 3056 6164 3064
rect 6140 3036 6148 3044
rect 6124 2936 6132 2944
rect 6236 3436 6244 3444
rect 6252 3316 6260 3324
rect 6220 3296 6228 3304
rect 6204 3276 6212 3284
rect 6252 3276 6260 3284
rect 6188 3236 6196 3244
rect 6220 3136 6228 3144
rect 6188 3096 6196 3104
rect 6204 3096 6212 3104
rect 6236 3116 6244 3124
rect 6220 3076 6228 3084
rect 6236 3036 6244 3044
rect 6172 3016 6180 3024
rect 6172 2996 6180 3004
rect 6284 3096 6292 3104
rect 6268 2996 6276 3004
rect 6252 2976 6260 2984
rect 6252 2956 6260 2964
rect 6268 2956 6276 2964
rect 6220 2936 6228 2944
rect 6140 2916 6148 2924
rect 6140 2896 6148 2904
rect 6108 2876 6116 2884
rect 6172 2916 6180 2924
rect 6204 2916 6212 2924
rect 6236 2916 6244 2924
rect 6156 2796 6164 2804
rect 6156 2776 6164 2784
rect 6124 2736 6132 2744
rect 6140 2736 6148 2744
rect 6156 2736 6164 2744
rect 6108 2696 6116 2704
rect 6124 2656 6132 2664
rect 6124 2596 6132 2604
rect 6124 2576 6132 2584
rect 6108 2536 6116 2544
rect 5980 2356 5988 2364
rect 6060 2356 6068 2364
rect 6044 2336 6052 2344
rect 5996 2276 6004 2284
rect 6012 2236 6020 2244
rect 6044 2256 6052 2264
rect 6108 2456 6116 2464
rect 6092 2436 6100 2444
rect 6028 2196 6036 2204
rect 6076 2196 6084 2204
rect 6092 2176 6100 2184
rect 6092 2156 6100 2164
rect 6076 2136 6084 2144
rect 6012 2116 6020 2124
rect 6060 2056 6068 2064
rect 6028 2016 6036 2024
rect 6044 2016 6052 2024
rect 5980 1956 5988 1964
rect 6012 1956 6020 1964
rect 5980 1916 5988 1924
rect 5996 1896 6004 1904
rect 6028 1896 6036 1904
rect 5964 1836 5972 1844
rect 5980 1796 5988 1804
rect 5980 1696 5988 1704
rect 5964 1636 5972 1644
rect 5980 1576 5988 1584
rect 5948 1536 5956 1544
rect 5948 1516 5952 1524
rect 5952 1516 5956 1524
rect 5932 1496 5940 1504
rect 5948 1496 5956 1504
rect 5916 1456 5924 1464
rect 5916 1416 5924 1424
rect 5900 1356 5908 1364
rect 5916 1296 5924 1304
rect 5900 1276 5908 1284
rect 5964 1416 5972 1424
rect 6028 1856 6036 1864
rect 6012 1836 6020 1844
rect 6012 1816 6020 1824
rect 6108 2076 6116 2084
rect 6092 2016 6100 2024
rect 6092 1956 6100 1964
rect 6060 1916 6068 1924
rect 6188 2796 6196 2804
rect 6236 2836 6244 2844
rect 6252 2816 6260 2824
rect 6156 2556 6164 2564
rect 6156 2536 6164 2544
rect 6156 2496 6164 2504
rect 6140 2376 6148 2384
rect 6156 2316 6164 2324
rect 6156 2276 6164 2284
rect 6140 2196 6148 2204
rect 6156 2076 6164 2084
rect 6156 2016 6164 2024
rect 6156 1976 6164 1984
rect 6156 1956 6164 1964
rect 6108 1936 6116 1944
rect 6124 1936 6132 1944
rect 6156 1936 6164 1944
rect 6108 1916 6116 1924
rect 6076 1876 6084 1884
rect 6076 1756 6084 1764
rect 6012 1536 6020 1544
rect 6044 1516 6052 1524
rect 6012 1496 6020 1504
rect 6028 1476 6036 1484
rect 5996 1376 6004 1384
rect 6044 1336 6052 1344
rect 6076 1496 6084 1504
rect 6140 1896 6148 1904
rect 6124 1876 6132 1884
rect 6108 1816 6116 1824
rect 6140 1716 6148 1724
rect 6108 1556 6116 1564
rect 6092 1476 6100 1484
rect 6092 1456 6100 1464
rect 6076 1376 6084 1384
rect 6012 1316 6020 1324
rect 6060 1316 6068 1324
rect 5980 1276 5988 1284
rect 5948 1236 5956 1244
rect 5932 1196 5940 1204
rect 5900 1176 5908 1184
rect 5884 1136 5892 1144
rect 5868 1116 5876 1124
rect 5884 1116 5892 1124
rect 5916 1136 5924 1144
rect 5868 1056 5876 1064
rect 5852 996 5860 1004
rect 5932 1076 5940 1084
rect 5836 956 5844 964
rect 5836 876 5844 884
rect 6028 1296 6036 1304
rect 5996 1236 6004 1244
rect 5964 1176 5972 1184
rect 6012 1196 6020 1204
rect 6012 1136 6020 1144
rect 6044 1136 6052 1144
rect 5980 1076 5988 1084
rect 5964 1056 5972 1064
rect 5996 1056 6004 1064
rect 5980 976 5988 984
rect 5996 976 6004 984
rect 5900 936 5908 944
rect 5916 936 5924 944
rect 5996 936 6004 944
rect 5884 876 5892 884
rect 5884 856 5892 864
rect 5852 816 5860 824
rect 5884 816 5892 824
rect 5836 756 5844 764
rect 5932 856 5940 864
rect 5980 816 5988 824
rect 6028 1056 6036 1064
rect 6044 1036 6052 1044
rect 6044 1016 6052 1024
rect 6028 976 6036 984
rect 6044 956 6052 964
rect 6028 876 6036 884
rect 6140 1616 6148 1624
rect 6124 1456 6132 1464
rect 6204 2696 6212 2704
rect 6188 2656 6196 2664
rect 6220 2656 6228 2664
rect 6188 2556 6196 2564
rect 6204 2516 6212 2524
rect 6220 2436 6228 2444
rect 6188 2376 6196 2384
rect 6268 2576 6276 2584
rect 6300 2596 6308 2604
rect 6268 2476 6276 2484
rect 6252 2356 6260 2364
rect 6204 2336 6212 2344
rect 6252 2336 6260 2344
rect 6188 2196 6196 2204
rect 6236 2256 6244 2264
rect 6220 2236 6228 2244
rect 6188 2016 6196 2024
rect 6188 1996 6196 2004
rect 6188 1956 6196 1964
rect 6204 1956 6212 1964
rect 6172 1876 6180 1884
rect 6204 1896 6212 1904
rect 6188 1856 6196 1864
rect 6156 1596 6164 1604
rect 6204 1816 6212 1824
rect 6188 1776 6196 1784
rect 6172 1476 6180 1484
rect 6108 1316 6116 1324
rect 6140 1276 6148 1284
rect 6124 1136 6132 1144
rect 6108 1116 6116 1124
rect 6076 1076 6084 1084
rect 6092 1076 6100 1084
rect 6076 1056 6084 1064
rect 6124 1076 6132 1084
rect 6108 1056 6116 1064
rect 6108 956 6116 964
rect 6076 896 6084 904
rect 6108 896 6116 904
rect 6060 876 6068 884
rect 6076 876 6084 884
rect 6044 816 6052 824
rect 6076 796 6084 804
rect 5916 776 5924 784
rect 5932 776 5940 784
rect 5788 696 5796 704
rect 5788 656 5796 664
rect 5740 596 5748 604
rect 5772 576 5780 584
rect 5708 536 5716 544
rect 5612 516 5620 524
rect 5628 516 5636 524
rect 5548 496 5556 504
rect 5596 476 5604 484
rect 5564 456 5572 464
rect 5580 456 5588 464
rect 5596 416 5604 424
rect 5484 396 5492 404
rect 5516 396 5524 404
rect 5468 356 5476 364
rect 5484 356 5492 364
rect 5532 356 5540 364
rect 5580 356 5588 364
rect 5404 336 5412 344
rect 5468 296 5476 304
rect 5436 276 5444 284
rect 5452 156 5460 164
rect 5532 316 5540 324
rect 5580 316 5588 324
rect 5644 456 5652 464
rect 5692 396 5700 404
rect 5708 396 5716 404
rect 5676 376 5684 384
rect 5660 316 5668 324
rect 5500 256 5508 264
rect 5516 256 5524 264
rect 5484 176 5492 184
rect 5500 176 5508 184
rect 5292 116 5300 124
rect 5260 76 5268 84
rect 5212 56 5220 64
rect 5228 56 5236 64
rect 5276 36 5284 44
rect 4908 16 4916 24
rect 5340 116 5348 124
rect 5388 136 5396 144
rect 5404 116 5412 124
rect 5468 76 5476 84
rect 5372 56 5380 64
rect 5532 156 5540 164
rect 5644 276 5652 284
rect 5740 476 5748 484
rect 5724 376 5732 384
rect 5724 336 5732 344
rect 5708 316 5716 324
rect 5580 196 5588 204
rect 5660 176 5668 184
rect 5564 96 5572 104
rect 5580 96 5588 104
rect 5628 96 5636 104
rect 5836 716 5844 724
rect 5820 696 5828 704
rect 5852 696 5860 704
rect 5900 756 5908 764
rect 5900 676 5908 684
rect 5884 656 5892 664
rect 5836 596 5844 604
rect 5868 596 5876 604
rect 5884 596 5892 604
rect 5804 576 5812 584
rect 5804 556 5812 564
rect 5788 476 5796 484
rect 5788 356 5796 364
rect 5788 336 5796 344
rect 5772 316 5780 324
rect 5804 276 5812 284
rect 5756 176 5764 184
rect 5708 136 5716 144
rect 5308 36 5316 44
rect 5676 56 5684 64
rect 5772 76 5780 84
rect 5916 636 5924 644
rect 6012 776 6020 784
rect 6092 756 6100 764
rect 6012 696 6020 704
rect 6076 696 6084 704
rect 6108 716 6116 724
rect 5948 656 5956 664
rect 5964 656 5972 664
rect 5996 656 6004 664
rect 6060 656 6068 664
rect 6092 656 6100 664
rect 5932 596 5940 604
rect 5948 576 5956 584
rect 5916 556 5924 564
rect 5932 556 5940 564
rect 5996 596 6004 604
rect 5852 536 5860 544
rect 5868 536 5876 544
rect 5964 536 5972 544
rect 5916 516 5924 524
rect 6060 556 6068 564
rect 6076 556 6084 564
rect 5964 496 5972 504
rect 5996 496 6004 504
rect 6012 496 6020 504
rect 5852 356 5860 364
rect 5932 336 5940 344
rect 5852 316 5860 324
rect 5884 316 5892 324
rect 5852 296 5860 304
rect 5948 296 5956 304
rect 5996 476 6004 484
rect 5980 396 5988 404
rect 5964 276 5972 284
rect 5836 196 5844 204
rect 5964 176 5972 184
rect 5932 136 5940 144
rect 6076 456 6084 464
rect 6028 396 6036 404
rect 6012 356 6020 364
rect 6012 336 6020 344
rect 6060 336 6068 344
rect 6060 296 6068 304
rect 5996 276 6004 284
rect 6028 256 6036 264
rect 6044 256 6052 264
rect 6044 216 6052 224
rect 6124 656 6132 664
rect 6124 636 6132 644
rect 6108 616 6116 624
rect 6252 2216 6260 2224
rect 6284 2316 6292 2324
rect 6268 2176 6276 2184
rect 6268 2076 6276 2084
rect 6300 1996 6308 2004
rect 6268 1956 6276 1964
rect 6252 1916 6260 1924
rect 6252 1896 6260 1904
rect 6236 1876 6244 1884
rect 6220 1796 6228 1804
rect 6220 1536 6228 1544
rect 6204 1496 6212 1504
rect 6204 1416 6212 1424
rect 6188 1376 6196 1384
rect 6188 1296 6196 1304
rect 6188 1276 6196 1284
rect 6188 1196 6196 1204
rect 6204 1196 6212 1204
rect 6172 1176 6180 1184
rect 6220 1176 6228 1184
rect 6188 1116 6196 1124
rect 6204 1116 6212 1124
rect 6220 1096 6228 1104
rect 6172 1076 6180 1084
rect 6188 1056 6196 1064
rect 6172 976 6180 984
rect 6268 1856 6276 1864
rect 6268 1596 6276 1604
rect 6268 1276 6276 1284
rect 6268 1256 6276 1264
rect 6252 1116 6260 1124
rect 6284 1076 6292 1084
rect 6268 1016 6276 1024
rect 6204 956 6212 964
rect 6236 956 6244 964
rect 6252 956 6260 964
rect 6156 736 6164 744
rect 6156 716 6164 724
rect 6236 936 6244 944
rect 6252 916 6260 924
rect 6252 876 6260 884
rect 6236 836 6244 844
rect 6252 756 6260 764
rect 6236 736 6244 744
rect 6140 576 6148 584
rect 6140 556 6148 564
rect 6156 556 6164 564
rect 6140 476 6148 484
rect 6092 436 6100 444
rect 6108 396 6116 404
rect 6092 356 6100 364
rect 6172 376 6180 384
rect 6252 716 6260 724
rect 6204 676 6212 684
rect 6220 676 6228 684
rect 6252 676 6260 684
rect 6220 616 6228 624
rect 6204 556 6212 564
rect 6204 476 6212 484
rect 6252 536 6260 544
rect 6284 916 6292 924
rect 6284 896 6292 904
rect 6284 836 6292 844
rect 6284 816 6292 824
rect 6284 736 6292 744
rect 6284 556 6292 564
rect 6284 516 6292 524
rect 6268 496 6276 504
rect 6220 416 6228 424
rect 6188 356 6196 364
rect 6140 316 6148 324
rect 6092 276 6100 284
rect 6124 276 6132 284
rect 6108 256 6116 264
rect 6076 216 6084 224
rect 6060 196 6068 204
rect 6156 236 6164 244
rect 6156 216 6164 224
rect 6252 256 6260 264
rect 6236 236 6244 244
rect 6204 196 6212 204
rect 6172 176 6180 184
rect 6236 176 6244 184
rect 6220 156 6228 164
rect 6268 156 6276 164
rect 6140 136 6148 144
rect 5964 116 5972 124
rect 6060 116 6068 124
rect 6124 116 6132 124
rect 5884 96 5892 104
rect 5900 96 5908 104
rect 5852 76 5860 84
rect 6028 56 6036 64
rect 5788 36 5796 44
rect 5468 16 5476 24
rect 5756 16 5764 24
<< metal3 >>
rect 1556 4617 1628 4623
rect 1732 4617 1756 4623
rect 1956 4617 1996 4623
rect 2420 4617 2460 4623
rect 2740 4617 2748 4623
rect 2900 4617 2908 4623
rect 3028 4617 3084 4623
rect 3476 4617 3500 4623
rect 3524 4617 4460 4623
rect 3112 4614 3160 4616
rect 3112 4606 3113 4614
rect 3122 4606 3123 4614
rect 3158 4606 3160 4614
rect 3112 4604 3160 4606
rect 404 4597 524 4603
rect 532 4597 2060 4603
rect 2132 4597 2924 4603
rect 2932 4597 3091 4603
rect 676 4577 732 4583
rect 740 4577 748 4583
rect 756 4577 1020 4583
rect 1028 4577 1068 4583
rect 1076 4577 2076 4583
rect 2292 4577 2396 4583
rect 3085 4583 3091 4597
rect 3220 4597 5196 4603
rect 5940 4597 6236 4603
rect 2868 4577 3075 4583
rect 3085 4577 3820 4583
rect 3069 4564 3075 4577
rect 4068 4577 4092 4583
rect 5844 4577 6172 4583
rect 980 4557 1260 4563
rect 1325 4557 2540 4563
rect 52 4537 108 4543
rect 116 4537 204 4543
rect 1325 4543 1331 4557
rect 2580 4557 2732 4563
rect 2932 4557 3052 4563
rect 3364 4557 3628 4563
rect 4708 4557 4812 4563
rect 4820 4557 4828 4563
rect 5364 4557 5596 4563
rect 5620 4557 5788 4563
rect 5940 4557 5996 4563
rect 6020 4557 6060 4563
rect 6100 4557 6156 4563
rect 1140 4537 1331 4543
rect 1380 4537 1580 4543
rect 1604 4537 1779 4543
rect -19 4517 12 4523
rect 100 4517 252 4523
rect 260 4517 460 4523
rect 484 4517 668 4523
rect 676 4517 716 4523
rect 868 4517 1100 4523
rect 1524 4517 1644 4523
rect 1684 4517 1740 4523
rect 1773 4523 1779 4537
rect 1796 4537 1804 4543
rect 2308 4537 2316 4543
rect 2452 4537 2684 4543
rect 2788 4537 2796 4543
rect 2964 4537 3260 4543
rect 3428 4537 3491 4543
rect 1773 4517 1916 4523
rect 2212 4517 2316 4523
rect 2676 4517 2700 4523
rect 2724 4517 2764 4523
rect 2772 4517 2780 4523
rect 2820 4517 2892 4523
rect 3069 4517 3164 4523
rect 628 4497 716 4503
rect 1028 4497 1084 4503
rect 1428 4497 1596 4503
rect 1636 4497 1740 4503
rect 1748 4497 1788 4503
rect 1908 4497 2044 4503
rect 2308 4497 2364 4503
rect 3069 4503 3075 4517
rect 3364 4517 3372 4523
rect 3380 4517 3420 4523
rect 3485 4523 3491 4537
rect 3508 4537 3516 4543
rect 4212 4537 4236 4543
rect 4244 4537 4716 4543
rect 4788 4537 4940 4543
rect 5444 4537 5484 4543
rect 5540 4537 5580 4543
rect 5588 4537 5740 4543
rect 5780 4537 5884 4543
rect 6004 4537 6156 4543
rect 3485 4517 3532 4523
rect 3972 4517 4140 4523
rect 4260 4517 4636 4523
rect 5268 4517 5324 4523
rect 5412 4517 5420 4523
rect 5469 4517 5548 4523
rect 3028 4497 3075 4503
rect 3092 4497 3484 4503
rect 3540 4497 3804 4503
rect 4148 4497 4204 4503
rect 4436 4497 4540 4503
rect 5108 4497 5324 4503
rect 5469 4503 5475 4517
rect 5556 4517 5692 4523
rect 5716 4517 5740 4523
rect 5764 4517 5788 4523
rect 5796 4517 5932 4523
rect 5428 4497 5475 4503
rect 5492 4497 5612 4503
rect 5684 4497 5756 4503
rect 5972 4497 6108 4503
rect 6164 4497 6172 4503
rect 6180 4497 6204 4503
rect 4141 4484 4147 4496
rect 1044 4477 1116 4483
rect 1348 4477 1660 4483
rect 1684 4477 1708 4483
rect 1940 4477 3020 4483
rect 3060 4477 3100 4483
rect 3380 4477 3660 4483
rect 4516 4477 4732 4483
rect 4740 4477 4780 4483
rect 5460 4477 5660 4483
rect 5988 4477 6012 4483
rect 372 4457 460 4463
rect 468 4457 732 4463
rect 740 4457 844 4463
rect 852 4457 1244 4463
rect 1252 4457 1276 4463
rect 1284 4457 1500 4463
rect 1517 4457 3052 4463
rect 1517 4443 1523 4457
rect 3124 4457 3452 4463
rect 3460 4457 3644 4463
rect 3908 4457 3948 4463
rect 3956 4457 4076 4463
rect 4084 4457 4348 4463
rect 4356 4457 4540 4463
rect 4548 4457 4572 4463
rect 4580 4457 4860 4463
rect 5060 4457 5244 4463
rect 5508 4457 5548 4463
rect 5556 4457 5580 4463
rect 5588 4457 5788 4463
rect 6164 4457 6284 4463
rect 1092 4437 1523 4443
rect 1620 4437 1644 4443
rect 2004 4437 2268 4443
rect 2285 4437 2332 4443
rect 2285 4423 2291 4437
rect 2388 4437 2396 4443
rect 2580 4437 4908 4443
rect 4916 4437 5020 4443
rect 5172 4437 5612 4443
rect 5636 4437 5740 4443
rect 6068 4437 6140 4443
rect 6148 4437 6188 4443
rect 1700 4417 2291 4423
rect 2308 4417 3644 4423
rect 3652 4417 4508 4423
rect 5156 4417 5884 4423
rect 6052 4417 6156 4423
rect 6164 4417 6236 4423
rect 1576 4414 1624 4416
rect 1576 4406 1577 4414
rect 1586 4406 1587 4414
rect 1622 4406 1624 4414
rect 1576 4404 1624 4406
rect 4664 4414 4712 4416
rect 4664 4406 4665 4414
rect 4674 4406 4675 4414
rect 4710 4406 4712 4414
rect 4664 4404 4712 4406
rect 1780 4397 3788 4403
rect 6004 4397 6028 4403
rect 1268 4377 1532 4383
rect 1556 4377 1580 4383
rect 1645 4377 1932 4383
rect 20 4357 236 4363
rect 1645 4363 1651 4377
rect 2100 4377 2284 4383
rect 2340 4377 2460 4383
rect 2660 4377 2732 4383
rect 2964 4377 5356 4383
rect 5380 4377 5388 4383
rect 5876 4377 6076 4383
rect 1524 4357 1651 4363
rect 1668 4357 1756 4363
rect 1780 4357 1900 4363
rect 1940 4357 2316 4363
rect 2324 4357 2684 4363
rect 2692 4357 2796 4363
rect 2804 4357 3596 4363
rect 3700 4357 3772 4363
rect 5236 4357 5468 4363
rect 5716 4357 5756 4363
rect 5764 4357 5820 4363
rect 5828 4357 5916 4363
rect 5956 4357 6028 4363
rect 6180 4357 6204 4363
rect 948 4337 1036 4343
rect 1492 4337 1740 4343
rect 1828 4337 2172 4343
rect 2180 4337 2556 4343
rect 2564 4337 2908 4343
rect 2916 4337 3276 4343
rect 3284 4337 3404 4343
rect 3412 4337 3500 4343
rect 3556 4337 3676 4343
rect 3684 4337 3692 4343
rect 5492 4337 5516 4343
rect 5796 4337 5852 4343
rect 5876 4337 5884 4343
rect 5892 4337 5916 4343
rect 6132 4337 6252 4343
rect 1540 4317 1788 4323
rect 2132 4317 2172 4323
rect 2244 4317 2284 4323
rect 2292 4317 2300 4323
rect 2388 4317 2428 4323
rect 2436 4317 2444 4323
rect 2836 4317 2924 4323
rect 2932 4317 2956 4323
rect 3188 4317 3372 4323
rect 3508 4317 3580 4323
rect 3620 4317 3884 4323
rect 4004 4317 4076 4323
rect 5108 4317 5164 4323
rect 5412 4317 5484 4323
rect 5524 4317 5580 4323
rect 5588 4317 5628 4323
rect 5908 4317 6220 4323
rect 1005 4304 1011 4316
rect 4205 4304 4211 4316
rect 148 4297 172 4303
rect 628 4297 828 4303
rect 1044 4297 1084 4303
rect 1204 4297 1772 4303
rect 1924 4297 1980 4303
rect 2308 4297 2524 4303
rect 2548 4297 2700 4303
rect 2756 4297 2844 4303
rect 2852 4297 2860 4303
rect 2884 4297 2940 4303
rect 2980 4297 3004 4303
rect 3012 4297 3020 4303
rect 3380 4297 3404 4303
rect 3412 4297 3436 4303
rect 3604 4297 3644 4303
rect 4276 4297 4284 4303
rect 4308 4297 4348 4303
rect 4356 4297 4444 4303
rect 4500 4297 4508 4303
rect 4516 4297 4556 4303
rect 4612 4297 4700 4303
rect 4916 4297 4956 4303
rect 4964 4297 5052 4303
rect 5076 4297 5180 4303
rect 5364 4297 5900 4303
rect 5908 4297 5932 4303
rect 3565 4284 3571 4296
rect 1284 4277 1372 4283
rect 1460 4277 1500 4283
rect 1508 4277 1964 4283
rect 2036 4277 2188 4283
rect 2212 4277 2316 4283
rect 2340 4277 2723 4283
rect 884 4257 988 4263
rect 1044 4257 1068 4263
rect 1124 4257 1404 4263
rect 1428 4257 1484 4263
rect 1540 4257 1580 4263
rect 1604 4257 1900 4263
rect 1988 4257 2700 4263
rect 2717 4263 2723 4277
rect 2861 4277 3212 4283
rect 2861 4263 2867 4277
rect 3236 4277 3420 4283
rect 3588 4277 3724 4283
rect 4084 4277 4092 4283
rect 4164 4277 4204 4283
rect 4276 4277 4300 4283
rect 4692 4277 4732 4283
rect 4740 4277 4748 4283
rect 5172 4277 5228 4283
rect 5380 4277 5420 4283
rect 5492 4277 5580 4283
rect 5604 4277 5660 4283
rect 5764 4277 5900 4283
rect 5940 4277 6172 4283
rect 6180 4277 6220 4283
rect 2717 4257 2867 4263
rect 2932 4257 2972 4263
rect 3060 4257 3500 4263
rect 3588 4257 3596 4263
rect 4132 4257 4188 4263
rect 4228 4257 4252 4263
rect 4660 4257 4860 4263
rect 5444 4257 5612 4263
rect 5620 4257 5692 4263
rect 5700 4257 5724 4263
rect 5748 4257 5788 4263
rect 5940 4257 5948 4263
rect 6036 4257 6044 4263
rect 6100 4257 6124 4263
rect 884 4237 1292 4243
rect 1332 4237 1356 4243
rect 1373 4237 1708 4243
rect 813 4224 819 4236
rect 829 4217 1100 4223
rect 212 4197 396 4203
rect 829 4203 835 4217
rect 1373 4223 1379 4237
rect 1812 4237 2508 4243
rect 2532 4237 2780 4243
rect 2788 4237 2924 4243
rect 2932 4237 3628 4243
rect 3652 4237 3996 4243
rect 4196 4237 4620 4243
rect 5396 4237 5676 4243
rect 5860 4237 5916 4243
rect 5924 4237 5980 4243
rect 1268 4217 1379 4223
rect 1396 4217 1468 4223
rect 1556 4217 2092 4223
rect 2868 4217 2924 4223
rect 3300 4217 3308 4223
rect 3412 4217 3420 4223
rect 3476 4217 3788 4223
rect 3988 4217 4076 4223
rect 4084 4217 4284 4223
rect 4596 4217 4604 4223
rect 5348 4217 5388 4223
rect 5469 4217 5500 4223
rect 3112 4214 3160 4216
rect 3112 4206 3113 4214
rect 3122 4206 3123 4214
rect 3158 4206 3160 4214
rect 3112 4204 3160 4206
rect 445 4197 835 4203
rect 196 4177 364 4183
rect 445 4183 451 4197
rect 868 4197 1052 4203
rect 1060 4197 2252 4203
rect 2388 4197 2908 4203
rect 2932 4197 2988 4203
rect 3236 4197 3347 4203
rect 388 4177 451 4183
rect 580 4177 652 4183
rect 669 4177 956 4183
rect 292 4157 332 4163
rect 372 4157 428 4163
rect 669 4163 675 4177
rect 980 4177 1628 4183
rect 1700 4177 1884 4183
rect 1924 4177 2028 4183
rect 2292 4177 2348 4183
rect 2388 4177 2492 4183
rect 2509 4177 3324 4183
rect 484 4157 675 4163
rect 708 4157 876 4163
rect 900 4157 972 4163
rect 1108 4157 1596 4163
rect 1620 4157 1660 4163
rect 1684 4157 1740 4163
rect 2509 4163 2515 4177
rect 3341 4183 3347 4197
rect 3444 4197 3628 4203
rect 3748 4197 3772 4203
rect 4084 4197 4227 4203
rect 3341 4177 3644 4183
rect 3764 4177 3964 4183
rect 3972 4177 4012 4183
rect 4020 4177 4204 4183
rect 4221 4183 4227 4197
rect 5252 4197 5420 4203
rect 5469 4203 5475 4217
rect 5812 4217 5868 4223
rect 5876 4217 5996 4223
rect 6196 4217 6220 4223
rect 5428 4197 5475 4203
rect 5860 4197 5916 4203
rect 5956 4197 6028 4203
rect 4221 4177 4396 4183
rect 5060 4177 5180 4183
rect 5188 4177 5276 4183
rect 5396 4177 5548 4183
rect 5556 4177 5660 4183
rect 5684 4177 6060 4183
rect 6132 4177 6156 4183
rect 1748 4157 2515 4163
rect 2644 4157 2828 4163
rect 2836 4157 3148 4163
rect 3156 4157 3308 4163
rect 3348 4157 3676 4163
rect 3700 4157 3715 4163
rect 132 4137 556 4143
rect 676 4137 684 4143
rect 692 4137 908 4143
rect 964 4137 1020 4143
rect 1044 4137 1356 4143
rect 1373 4137 1420 4143
rect 148 4117 188 4123
rect 212 4117 412 4123
rect 756 4117 931 4123
rect 356 4097 396 4103
rect 612 4097 636 4103
rect 925 4103 931 4117
rect 996 4117 1004 4123
rect 1012 4117 1036 4123
rect 1092 4117 1228 4123
rect 1252 4117 1260 4123
rect 1373 4123 1379 4137
rect 1444 4137 1500 4143
rect 1508 4137 2812 4143
rect 2845 4137 3036 4143
rect 1348 4117 1379 4123
rect 1796 4117 1932 4123
rect 1940 4117 1964 4123
rect 1972 4117 1980 4123
rect 2068 4117 2284 4123
rect 2292 4117 2412 4123
rect 2452 4117 2556 4123
rect 2564 4117 2668 4123
rect 2845 4123 2851 4137
rect 3044 4137 3276 4143
rect 3348 4137 3404 4143
rect 3620 4137 3692 4143
rect 3709 4143 3715 4157
rect 3732 4157 4172 4163
rect 4372 4157 4380 4163
rect 5044 4157 5084 4163
rect 5092 4157 5116 4163
rect 5268 4157 5468 4163
rect 5940 4157 5980 4163
rect 6068 4157 6124 4163
rect 3709 4137 3820 4143
rect 3940 4137 4028 4143
rect 4052 4137 4115 4143
rect 2676 4117 2851 4123
rect 2868 4117 2940 4123
rect 2948 4117 3004 4123
rect 3028 4117 3084 4123
rect 3252 4117 3340 4123
rect 3364 4117 3468 4123
rect 3572 4117 3612 4123
rect 3668 4117 3980 4123
rect 4036 4117 4092 4123
rect 4109 4123 4115 4137
rect 4212 4137 4236 4143
rect 4244 4137 4300 4143
rect 4324 4137 4716 4143
rect 4724 4137 4780 4143
rect 5101 4137 5244 4143
rect 5101 4124 5107 4137
rect 5268 4137 5404 4143
rect 5412 4137 5564 4143
rect 5684 4137 5692 4143
rect 5700 4137 5740 4143
rect 5796 4137 6044 4143
rect 6052 4137 6268 4143
rect 4109 4117 4204 4123
rect 4244 4117 4300 4123
rect 4308 4117 4364 4123
rect 4596 4117 4764 4123
rect 4964 4117 5020 4123
rect 5252 4117 5292 4123
rect 5300 4117 5324 4123
rect 5380 4117 5436 4123
rect 5492 4117 5548 4123
rect 5716 4117 5772 4123
rect 5892 4117 5900 4123
rect 5908 4117 6028 4123
rect 6180 4117 6220 4123
rect 925 4097 988 4103
rect 1012 4097 1308 4103
rect 1316 4097 1356 4103
rect 1364 4097 1468 4103
rect 1476 4097 1548 4103
rect 1556 4097 1644 4103
rect 1684 4097 1740 4103
rect 1876 4097 1964 4103
rect 1988 4097 2156 4103
rect 2196 4097 2380 4103
rect 2404 4097 2492 4103
rect 2516 4097 2524 4103
rect 2548 4097 2604 4103
rect 2628 4097 3020 4103
rect 3076 4097 3196 4103
rect 3236 4097 3308 4103
rect 3620 4097 3708 4103
rect 3716 4097 3836 4103
rect 3844 4097 3916 4103
rect 4180 4097 4332 4103
rect 4388 4097 4396 4103
rect 4756 4097 4940 4103
rect 5156 4097 5164 4103
rect 5236 4097 5292 4103
rect 5332 4097 5356 4103
rect 5684 4097 5740 4103
rect 5748 4097 5916 4103
rect 5924 4097 6188 4103
rect 6228 4097 6284 4103
rect 205 4084 211 4096
rect 324 4077 364 4083
rect 468 4077 876 4083
rect 932 4077 988 4083
rect 1028 4077 1100 4083
rect 1780 4077 1836 4083
rect 1876 4077 2220 4083
rect 2420 4077 2572 4083
rect 2596 4077 2668 4083
rect 2724 4077 2780 4083
rect 2788 4077 2812 4083
rect 2820 4077 2876 4083
rect 2916 4077 2972 4083
rect 2980 4077 3100 4083
rect 3268 4077 3276 4083
rect 3380 4077 3468 4083
rect 3572 4077 3660 4083
rect 3668 4077 3724 4083
rect 3732 4077 3852 4083
rect 3860 4077 3900 4083
rect 3988 4077 4076 4083
rect 4100 4077 4268 4083
rect 5876 4077 5932 4083
rect 6036 4077 6060 4083
rect 6132 4077 6284 4083
rect 84 4057 364 4063
rect 916 4057 972 4063
rect 980 4057 1084 4063
rect 1092 4057 1148 4063
rect 1156 4057 1212 4063
rect 1236 4057 1324 4063
rect 1396 4057 1532 4063
rect 1556 4057 1692 4063
rect 1700 4057 1756 4063
rect 1828 4057 1852 4063
rect 1892 4057 1900 4063
rect 1908 4057 1932 4063
rect 1940 4057 1971 4063
rect 996 4037 1116 4043
rect 1300 4037 1516 4043
rect 1524 4037 1692 4043
rect 1716 4037 1788 4043
rect 1844 4037 1948 4043
rect 1965 4043 1971 4057
rect 2004 4057 2860 4063
rect 2868 4057 2988 4063
rect 2996 4057 3388 4063
rect 3396 4057 3596 4063
rect 3604 4057 4236 4063
rect 4244 4057 4268 4063
rect 4276 4057 4556 4063
rect 4564 4057 4700 4063
rect 5220 4057 5420 4063
rect 5428 4057 5484 4063
rect 5844 4057 6060 4063
rect 1965 4037 2124 4043
rect 2308 4037 2316 4043
rect 2388 4037 2556 4043
rect 2580 4037 5980 4043
rect 5997 4037 6115 4043
rect 884 4017 1196 4023
rect 1236 4017 1340 4023
rect 1460 4017 1484 4023
rect 1492 4017 1516 4023
rect 1668 4017 1980 4023
rect 2036 4017 2092 4023
rect 2164 4017 2444 4023
rect 2452 4017 2636 4023
rect 2836 4017 4620 4023
rect 5188 4017 5228 4023
rect 5364 4017 5756 4023
rect 5764 4017 5852 4023
rect 5997 4023 6003 4037
rect 5956 4017 6003 4023
rect 6109 4023 6115 4037
rect 6132 4037 6220 4043
rect 6109 4017 6140 4023
rect 1576 4014 1624 4016
rect 1576 4006 1577 4014
rect 1586 4006 1587 4014
rect 1622 4006 1624 4014
rect 1576 4004 1624 4006
rect 4664 4014 4712 4016
rect 4664 4006 4665 4014
rect 4674 4006 4675 4014
rect 4710 4006 4712 4014
rect 4664 4004 4712 4006
rect 788 3997 940 4003
rect 948 3997 1292 4003
rect 1396 3997 1436 4003
rect 1460 3997 1516 4003
rect 2084 3997 2540 4003
rect 2564 3997 2668 4003
rect 2740 3997 2764 4003
rect 2868 3997 2876 4003
rect 2900 3997 3532 4003
rect 3556 3997 3596 4003
rect 3604 3997 3612 4003
rect 3652 3997 3660 4003
rect 3700 3997 3884 4003
rect 3908 3997 4012 4003
rect 4052 3997 4172 4003
rect 4228 3997 4284 4003
rect 4292 3997 4348 4003
rect 4436 3997 4460 4003
rect 4468 3997 4636 4003
rect 5380 3997 5788 4003
rect 5860 3997 5884 4003
rect 5972 3997 6156 4003
rect 1044 3977 1116 3983
rect 1140 3977 1180 3983
rect 1204 3977 1388 3983
rect 1396 3977 1452 3983
rect 1700 3977 1756 3983
rect 1773 3977 1868 3983
rect 84 3957 268 3963
rect 276 3957 284 3963
rect 1076 3957 1132 3963
rect 1773 3963 1779 3977
rect 1908 3977 2028 3983
rect 2068 3977 2444 3983
rect 2468 3977 2604 3983
rect 2660 3977 2748 3983
rect 2772 3977 2796 3983
rect 2804 3977 3372 3983
rect 3380 3977 4140 3983
rect 4148 3977 4284 3983
rect 4292 3977 4348 3983
rect 4356 3977 4588 3983
rect 4596 3977 4780 3983
rect 5908 3977 5996 3983
rect 6036 3977 6060 3983
rect 1172 3957 1779 3963
rect 2212 3957 2476 3963
rect 2500 3957 2860 3963
rect 2884 3957 3564 3963
rect 3572 3957 3948 3963
rect 3956 3957 4012 3963
rect 4020 3957 4364 3963
rect 5796 3957 5932 3963
rect 6020 3957 6076 3963
rect 260 3937 332 3943
rect 900 3937 1404 3943
rect 1460 3937 2028 3943
rect 2388 3937 2428 3943
rect 2452 3937 2636 3943
rect 2724 3937 2780 3943
rect 2788 3937 2956 3943
rect 2964 3937 3116 3943
rect 3124 3937 3420 3943
rect 3444 3940 3532 3943
rect 3437 3937 3532 3940
rect 3588 3937 3596 3943
rect 4068 3937 4076 3943
rect 4148 3937 4156 3943
rect 4212 3937 4236 3943
rect 5060 3937 5084 3943
rect 5396 3937 5740 3943
rect 5780 3937 5884 3943
rect 5908 3937 5932 3943
rect 6004 3937 6284 3943
rect 100 3917 204 3923
rect 317 3917 332 3923
rect 84 3897 124 3903
rect 180 3897 275 3903
rect 116 3877 156 3883
rect 180 3877 204 3883
rect 244 3877 252 3883
rect 269 3883 275 3897
rect 317 3903 323 3917
rect 340 3917 412 3923
rect 692 3917 860 3923
rect 1028 3917 1148 3923
rect 1188 3917 1228 3923
rect 1252 3917 1260 3923
rect 1492 3917 1868 3923
rect 2004 3917 2012 3923
rect 2068 3917 2140 3923
rect 2164 3917 2252 3923
rect 2340 3917 2492 3923
rect 2548 3917 2636 3923
rect 2676 3917 2732 3923
rect 2772 3917 2780 3923
rect 2868 3917 3340 3923
rect 3380 3917 3404 3923
rect 3437 3920 3452 3923
rect 3444 3917 3452 3920
rect 3476 3917 3740 3923
rect 3949 3923 3955 3936
rect 3748 3917 3980 3923
rect 3988 3917 4060 3923
rect 4116 3917 4124 3923
rect 4180 3917 4220 3923
rect 4276 3917 4460 3923
rect 4996 3917 5068 3923
rect 5204 3917 5228 3923
rect 5236 3917 5244 3923
rect 5332 3917 5404 3923
rect 5444 3917 5580 3923
rect 5588 3917 5676 3923
rect 5844 3917 5948 3923
rect 5988 3917 6124 3923
rect 6164 3917 6220 3923
rect 292 3897 323 3903
rect 356 3897 412 3903
rect 420 3897 556 3903
rect 868 3897 908 3903
rect 1012 3897 1084 3903
rect 1213 3897 1571 3903
rect 269 3877 460 3883
rect 532 3877 572 3883
rect 580 3877 636 3883
rect 852 3877 1068 3883
rect 1213 3883 1219 3897
rect 1092 3877 1219 3883
rect 1364 3877 1427 3883
rect 148 3857 156 3863
rect 212 3857 220 3863
rect 228 3857 508 3863
rect 964 3857 972 3863
rect 1076 3857 1084 3863
rect 1140 3857 1196 3863
rect 1421 3863 1427 3877
rect 1444 3877 1548 3883
rect 1565 3883 1571 3897
rect 1604 3897 2060 3903
rect 2388 3897 2396 3903
rect 2436 3897 2892 3903
rect 2996 3897 3212 3903
rect 3268 3897 3308 3903
rect 3412 3897 3500 3903
rect 3668 3897 3676 3903
rect 3700 3897 3740 3903
rect 3860 3897 4252 3903
rect 4077 3884 4083 3897
rect 4356 3897 4508 3903
rect 4772 3897 4963 3903
rect 1565 3877 1804 3883
rect 1828 3877 1836 3883
rect 1908 3877 1964 3883
rect 2004 3877 2108 3883
rect 2148 3877 2396 3883
rect 2436 3877 2476 3883
rect 2596 3877 2620 3883
rect 2660 3877 2668 3883
rect 2756 3877 2780 3883
rect 2820 3877 2860 3883
rect 2916 3877 3020 3883
rect 3028 3877 3468 3883
rect 3476 3877 3548 3883
rect 3572 3877 3692 3883
rect 3732 3877 4060 3883
rect 4100 3877 4284 3883
rect 4564 3877 4796 3883
rect 4804 3877 4940 3883
rect 4957 3883 4963 3897
rect 5060 3897 5091 3903
rect 4957 3877 5052 3883
rect 5085 3883 5091 3897
rect 5172 3897 5260 3903
rect 5348 3897 5452 3903
rect 5476 3897 5596 3903
rect 5604 3897 5660 3903
rect 5668 3897 5708 3903
rect 5748 3897 5772 3903
rect 5780 3897 5820 3903
rect 5876 3897 5916 3903
rect 6116 3897 6124 3903
rect 6132 3897 6188 3903
rect 5085 3877 5100 3883
rect 5124 3877 5196 3883
rect 5252 3877 5292 3883
rect 5412 3877 5772 3883
rect 5780 3877 5836 3883
rect 6004 3877 6028 3883
rect 6068 3877 6124 3883
rect 6132 3877 6188 3883
rect 1268 3857 1411 3863
rect 1421 3857 1484 3863
rect 148 3837 236 3843
rect 324 3837 364 3843
rect 388 3837 508 3843
rect 516 3837 908 3843
rect 1012 3837 1164 3843
rect 1204 3837 1228 3843
rect 1268 3837 1340 3843
rect 1405 3843 1411 3857
rect 1524 3857 1564 3863
rect 1780 3857 2019 3863
rect 1405 3837 1436 3843
rect 1460 3837 1612 3843
rect 1716 3837 1740 3843
rect 1812 3837 1980 3843
rect 2013 3843 2019 3857
rect 2068 3857 2092 3863
rect 2164 3857 2188 3863
rect 2196 3857 2412 3863
rect 2452 3857 2524 3863
rect 2564 3857 2604 3863
rect 2692 3857 2716 3863
rect 2724 3857 2828 3863
rect 2836 3857 2892 3863
rect 2900 3857 3756 3863
rect 3764 3857 3948 3863
rect 3956 3857 4140 3863
rect 4164 3857 4188 3863
rect 5188 3857 5244 3863
rect 5252 3857 5356 3863
rect 5540 3857 5628 3863
rect 5716 3857 5836 3863
rect 5844 3857 5868 3863
rect 5924 3857 5964 3863
rect 5972 3857 6140 3863
rect 6164 3857 6204 3863
rect 2013 3837 2060 3843
rect 2116 3837 2243 3843
rect 260 3817 636 3823
rect 820 3817 1500 3823
rect 1508 3817 2028 3823
rect 2036 3817 2220 3823
rect 2237 3823 2243 3837
rect 2292 3837 2348 3843
rect 2404 3837 3212 3843
rect 3252 3837 3260 3843
rect 3316 3837 3324 3843
rect 3348 3837 3596 3843
rect 3636 3837 3692 3843
rect 4004 3837 4396 3843
rect 5364 3837 5788 3843
rect 5908 3837 6028 3843
rect 6164 3837 6284 3843
rect 2237 3817 3068 3823
rect 3412 3817 4588 3823
rect 4596 3817 4620 3823
rect 4708 3817 4972 3823
rect 5268 3817 5292 3823
rect 5428 3817 5676 3823
rect 5684 3817 5836 3823
rect 6020 3817 6044 3823
rect 6164 3817 6172 3823
rect 3112 3814 3160 3816
rect 3112 3806 3113 3814
rect 3122 3806 3123 3814
rect 3158 3806 3160 3814
rect 3112 3804 3160 3806
rect 244 3797 268 3803
rect 276 3797 332 3803
rect 404 3797 460 3803
rect 484 3797 700 3803
rect 820 3797 940 3803
rect 948 3797 1411 3803
rect 29 3777 44 3783
rect 29 3743 35 3777
rect 100 3777 124 3783
rect 212 3777 284 3783
rect 308 3777 588 3783
rect 596 3777 844 3783
rect 852 3777 1116 3783
rect 1124 3777 1276 3783
rect 1405 3783 1411 3797
rect 1428 3797 1708 3803
rect 1748 3797 1795 3803
rect 1405 3777 1708 3783
rect 1748 3780 1772 3783
rect 1789 3783 1795 3797
rect 1892 3797 1916 3803
rect 1988 3797 2220 3803
rect 2372 3797 2604 3803
rect 2644 3797 2860 3803
rect 2868 3797 2924 3803
rect 3060 3797 3084 3803
rect 3188 3797 3772 3803
rect 3892 3797 3980 3803
rect 4004 3797 4156 3803
rect 4196 3797 5084 3803
rect 5092 3797 5132 3803
rect 5204 3797 5276 3803
rect 5748 3797 5804 3803
rect 6004 3797 6156 3803
rect 6196 3797 6220 3803
rect 1748 3777 1779 3780
rect 1789 3777 2076 3783
rect 2196 3777 2508 3783
rect 2548 3777 2668 3783
rect 2692 3777 3324 3783
rect 3540 3777 3795 3783
rect 3789 3764 3795 3777
rect 3821 3777 4252 3783
rect 3821 3764 3827 3777
rect 4276 3777 5660 3783
rect 5668 3777 5676 3783
rect 5684 3777 5804 3783
rect 5828 3777 5836 3783
rect 6052 3777 6060 3783
rect 6100 3777 6124 3783
rect 308 3757 524 3763
rect 916 3757 1084 3763
rect 1108 3757 1132 3763
rect 1204 3757 1420 3763
rect 1444 3757 1468 3763
rect 1524 3757 1660 3763
rect 1773 3760 1900 3763
rect 1780 3757 1900 3760
rect 1924 3757 2748 3763
rect 2820 3757 2908 3763
rect 2932 3757 3020 3763
rect 3060 3757 3180 3763
rect 3188 3757 3308 3763
rect 3316 3757 3372 3763
rect 3476 3757 3532 3763
rect 3645 3757 3676 3763
rect 29 3737 51 3743
rect 45 3723 51 3737
rect 68 3737 92 3743
rect 132 3737 140 3743
rect 212 3737 316 3743
rect 372 3737 396 3743
rect 468 3737 476 3743
rect 500 3737 540 3743
rect 836 3737 860 3743
rect 932 3737 956 3743
rect 1076 3737 1116 3743
rect 1140 3737 1148 3743
rect 1156 3737 1372 3743
rect 1437 3737 1468 3743
rect 1389 3724 1395 3736
rect 45 3717 76 3723
rect 100 3717 124 3723
rect 148 3717 268 3723
rect 372 3717 396 3723
rect 420 3717 540 3723
rect 548 3717 620 3723
rect 820 3717 876 3723
rect 1012 3717 1148 3723
rect 1156 3717 1228 3723
rect 148 3697 204 3703
rect 244 3697 524 3703
rect 548 3697 556 3703
rect 564 3697 588 3703
rect 644 3697 668 3703
rect 916 3697 1052 3703
rect 1076 3697 1116 3703
rect 1140 3697 1244 3703
rect 1268 3697 1404 3703
rect 1437 3703 1443 3737
rect 1492 3737 1564 3743
rect 1620 3737 1724 3743
rect 1860 3737 1884 3743
rect 1892 3737 1932 3743
rect 2020 3737 2348 3743
rect 2372 3737 2444 3743
rect 2548 3737 2684 3743
rect 2708 3737 2828 3743
rect 2893 3737 3315 3743
rect 1460 3717 1468 3723
rect 1492 3717 1516 3723
rect 1556 3717 1651 3723
rect 1437 3697 1475 3703
rect 404 3677 556 3683
rect 948 3677 988 3683
rect 996 3677 1100 3683
rect 1108 3677 1164 3683
rect 1188 3677 1452 3683
rect 1469 3683 1475 3697
rect 1492 3697 1612 3703
rect 1645 3703 1651 3717
rect 1668 3717 1676 3723
rect 1684 3717 1779 3723
rect 1645 3697 1676 3703
rect 1732 3697 1740 3703
rect 1773 3703 1779 3717
rect 1812 3717 2028 3723
rect 2068 3717 2108 3723
rect 2164 3717 2252 3723
rect 2324 3717 2444 3723
rect 2461 3723 2467 3736
rect 2461 3717 2636 3723
rect 2676 3717 2764 3723
rect 2788 3717 2860 3723
rect 2893 3723 2899 3737
rect 3309 3724 3315 3737
rect 3524 3737 3580 3743
rect 3620 3737 3628 3743
rect 2884 3717 2899 3723
rect 2916 3717 3260 3723
rect 3284 3717 3292 3723
rect 3396 3717 3420 3723
rect 3645 3723 3651 3757
rect 3732 3757 3772 3763
rect 3828 3757 3852 3763
rect 3972 3757 4012 3763
rect 4100 3757 4556 3763
rect 5252 3757 5372 3763
rect 5444 3757 5484 3763
rect 5524 3757 5548 3763
rect 5732 3757 5900 3763
rect 6237 3757 6284 3763
rect 3812 3737 3820 3743
rect 3828 3737 3868 3743
rect 3876 3737 4108 3743
rect 4116 3737 4172 3743
rect 4189 3737 4236 3743
rect 3524 3717 3651 3723
rect 3668 3717 3763 3723
rect 1773 3697 1852 3703
rect 1876 3697 1916 3703
rect 1972 3697 2092 3703
rect 2116 3697 2188 3703
rect 2292 3697 2412 3703
rect 2468 3697 2508 3703
rect 2516 3697 2604 3703
rect 2676 3697 2700 3703
rect 2740 3697 2828 3703
rect 3012 3697 3020 3703
rect 3044 3697 3155 3703
rect 1469 3677 1484 3683
rect 1604 3677 1708 3683
rect 1748 3677 1884 3683
rect 1892 3677 2252 3683
rect 2388 3677 2428 3683
rect 2452 3677 2492 3683
rect 2516 3677 2700 3683
rect 2740 3677 2892 3683
rect 2916 3677 2956 3683
rect 2980 3677 3068 3683
rect 3092 3677 3132 3683
rect 3149 3683 3155 3697
rect 3236 3697 3612 3703
rect 3636 3697 3740 3703
rect 3757 3703 3763 3717
rect 3796 3717 3948 3723
rect 4052 3717 4140 3723
rect 4189 3723 4195 3737
rect 4244 3737 4300 3743
rect 4564 3737 4636 3743
rect 4884 3737 4940 3743
rect 5188 3737 5324 3743
rect 5396 3737 5452 3743
rect 5476 3737 5644 3743
rect 5652 3737 5964 3743
rect 6237 3743 6243 3757
rect 6036 3737 6243 3743
rect 6260 3737 6284 3743
rect 4164 3717 4195 3723
rect 4228 3717 4236 3723
rect 4292 3717 4460 3723
rect 4548 3717 4556 3723
rect 4596 3717 4604 3723
rect 5044 3717 5148 3723
rect 5236 3717 5372 3723
rect 5444 3717 5516 3723
rect 5540 3717 5580 3723
rect 5636 3717 5724 3723
rect 5732 3717 5740 3723
rect 5796 3717 5884 3723
rect 5908 3717 5932 3723
rect 6052 3717 6140 3723
rect 3981 3704 3987 3716
rect 3757 3697 3820 3703
rect 4020 3697 4060 3703
rect 4068 3697 4124 3703
rect 4596 3697 4828 3703
rect 5012 3697 5116 3703
rect 5156 3697 5292 3703
rect 5332 3697 5356 3703
rect 5380 3697 5708 3703
rect 5732 3697 5756 3703
rect 5844 3697 5884 3703
rect 6036 3697 6124 3703
rect 6132 3697 6172 3703
rect 6196 3697 6204 3703
rect 6212 3697 6236 3703
rect 6260 3697 6284 3703
rect 3149 3677 3244 3683
rect 3268 3677 3475 3683
rect 308 3657 428 3663
rect 468 3657 908 3663
rect 1044 3657 1580 3663
rect 1620 3657 2108 3663
rect 2180 3657 2332 3663
rect 2356 3657 2716 3663
rect 2772 3657 2828 3663
rect 2868 3657 2972 3663
rect 3012 3657 3148 3663
rect 3284 3657 3324 3663
rect 3348 3657 3404 3663
rect 3412 3657 3436 3663
rect 3469 3663 3475 3677
rect 3492 3677 3836 3683
rect 3860 3677 3980 3683
rect 4084 3677 4188 3683
rect 4260 3677 4396 3683
rect 4628 3677 5468 3683
rect 5620 3677 5676 3683
rect 5732 3677 5820 3683
rect 6116 3677 6124 3683
rect 3469 3657 5484 3663
rect 5556 3657 5756 3663
rect 5780 3657 5900 3663
rect 973 3644 979 3656
rect 36 3637 140 3643
rect 148 3637 332 3643
rect 340 3637 428 3643
rect 436 3637 620 3643
rect 1044 3637 1836 3643
rect 1844 3637 2604 3643
rect 2612 3637 3596 3643
rect 3620 3637 5084 3643
rect 5092 3637 5164 3643
rect 5188 3637 5324 3643
rect 5332 3637 5452 3643
rect 5460 3637 5516 3643
rect 5524 3637 5836 3643
rect 5844 3637 5916 3643
rect 5924 3637 6012 3643
rect 244 3617 604 3623
rect 612 3617 1036 3623
rect 1060 3617 1180 3623
rect 1396 3617 1532 3623
rect 1684 3617 1900 3623
rect 1908 3617 2012 3623
rect 2036 3617 2060 3623
rect 2068 3617 2300 3623
rect 2308 3617 2476 3623
rect 2676 3617 2780 3623
rect 2836 3617 2908 3623
rect 3076 3617 3116 3623
rect 3188 3617 3372 3623
rect 3396 3617 3420 3623
rect 3428 3617 3436 3623
rect 3460 3617 3660 3623
rect 3668 3617 3932 3623
rect 3940 3617 4172 3623
rect 4180 3617 4236 3623
rect 4388 3617 4636 3623
rect 5332 3617 5356 3623
rect 5508 3617 5564 3623
rect 5604 3617 5836 3623
rect 5844 3617 5852 3623
rect 5940 3617 5964 3623
rect 5988 3617 6028 3623
rect 1576 3614 1624 3616
rect 1576 3606 1577 3614
rect 1586 3606 1587 3614
rect 1622 3606 1624 3614
rect 1576 3604 1624 3606
rect 4664 3614 4712 3616
rect 4664 3606 4665 3614
rect 4674 3606 4675 3614
rect 4710 3606 4712 3614
rect 4664 3604 4712 3606
rect 52 3597 76 3603
rect 132 3597 140 3603
rect 212 3597 492 3603
rect 660 3597 748 3603
rect 772 3597 876 3603
rect 1069 3597 1084 3603
rect 580 3577 636 3583
rect 1069 3583 1075 3597
rect 1140 3597 1331 3603
rect 820 3577 1075 3583
rect 1092 3577 1132 3583
rect 1172 3577 1212 3583
rect 1325 3583 1331 3597
rect 1348 3597 1468 3603
rect 1844 3597 1868 3603
rect 2116 3597 2236 3603
rect 2468 3597 2508 3603
rect 2564 3597 2572 3603
rect 2580 3597 2700 3603
rect 2724 3597 2764 3603
rect 2804 3597 2860 3603
rect 2980 3597 3052 3603
rect 3076 3597 3180 3603
rect 3332 3597 3820 3603
rect 3844 3597 4028 3603
rect 4036 3597 4044 3603
rect 4068 3597 4588 3603
rect 5316 3597 5788 3603
rect 1325 3577 1612 3583
rect 1700 3577 1836 3583
rect 1860 3577 2204 3583
rect 2228 3577 2380 3583
rect 2420 3577 2524 3583
rect 3092 3577 5196 3583
rect 5204 3577 5276 3583
rect 5332 3577 5420 3583
rect 5533 3577 5852 3583
rect 84 3557 204 3563
rect 356 3557 844 3563
rect 964 3557 1052 3563
rect 1124 3557 1180 3563
rect 1364 3557 1436 3563
rect 1444 3557 1619 3563
rect 276 3537 284 3543
rect 564 3537 764 3543
rect 804 3537 860 3543
rect 900 3537 1004 3543
rect 1124 3537 1228 3543
rect 1316 3537 1372 3543
rect 1380 3537 1484 3543
rect 1565 3537 1596 3543
rect 557 3524 563 3536
rect 68 3517 204 3523
rect 404 3517 412 3523
rect 596 3517 604 3523
rect 660 3517 700 3523
rect 900 3517 908 3523
rect 980 3517 1116 3523
rect 1124 3517 1148 3523
rect 1188 3517 1244 3523
rect 1268 3517 1292 3523
rect 1332 3517 1340 3523
rect 1364 3517 1388 3523
rect 1565 3523 1571 3537
rect 1613 3543 1619 3557
rect 1636 3557 1692 3563
rect 1716 3557 1900 3563
rect 1956 3557 2028 3563
rect 2036 3557 2092 3563
rect 2100 3557 2156 3563
rect 2164 3557 2435 3563
rect 2429 3544 2435 3557
rect 2452 3557 2540 3563
rect 2612 3557 2732 3563
rect 2836 3557 2876 3563
rect 3028 3557 3100 3563
rect 3220 3557 3244 3563
rect 3316 3557 3356 3563
rect 3476 3557 3532 3563
rect 3572 3557 3724 3563
rect 3732 3557 3756 3563
rect 3828 3557 3964 3563
rect 3988 3557 4012 3563
rect 4020 3557 4060 3563
rect 4100 3557 4236 3563
rect 4260 3557 4380 3563
rect 5533 3563 5539 3577
rect 5956 3577 5980 3583
rect 4596 3557 5539 3563
rect 5556 3557 6076 3563
rect 5901 3544 5907 3557
rect 6084 3557 6140 3563
rect 1613 3537 1692 3543
rect 1780 3537 1884 3543
rect 1924 3537 1964 3543
rect 2036 3537 2316 3543
rect 2340 3537 2396 3543
rect 2452 3537 2620 3543
rect 2660 3537 2796 3543
rect 2852 3537 3212 3543
rect 3236 3537 3292 3543
rect 3316 3537 3916 3543
rect 3924 3537 4172 3543
rect 4212 3537 4732 3543
rect 5236 3537 5244 3543
rect 5316 3537 5500 3543
rect 5757 3537 5772 3543
rect 1540 3517 1571 3523
rect 1940 3517 2003 3523
rect 52 3497 76 3503
rect 132 3497 172 3503
rect 180 3497 268 3503
rect 276 3497 316 3503
rect 573 3503 579 3516
rect 404 3497 579 3503
rect 612 3497 636 3503
rect 692 3497 812 3503
rect 820 3497 1260 3503
rect 1284 3497 1404 3503
rect 1412 3497 1516 3503
rect 1540 3497 1580 3503
rect 1597 3497 1660 3503
rect 52 3477 188 3483
rect 228 3477 348 3483
rect 404 3477 428 3483
rect 500 3477 540 3483
rect 580 3477 604 3483
rect 612 3477 620 3483
rect 628 3477 780 3483
rect 804 3477 844 3483
rect 868 3477 892 3483
rect 980 3477 1020 3483
rect 1108 3477 1196 3483
rect 1300 3477 1356 3483
rect 1380 3477 1436 3483
rect 1597 3483 1603 3497
rect 1700 3497 1804 3503
rect 1997 3503 2003 3517
rect 2020 3517 2044 3523
rect 2084 3517 2348 3523
rect 2388 3517 2531 3523
rect 1997 3497 2019 3503
rect 1492 3477 1603 3483
rect 1620 3477 1708 3483
rect 1780 3477 1868 3483
rect 2013 3483 2019 3497
rect 2084 3497 2188 3503
rect 2212 3497 2412 3503
rect 2436 3497 2460 3503
rect 2525 3503 2531 3517
rect 2564 3517 2892 3523
rect 2948 3517 2988 3523
rect 3700 3517 3900 3523
rect 3924 3517 3964 3523
rect 3988 3517 4108 3523
rect 4244 3517 4316 3523
rect 4468 3517 4556 3523
rect 4564 3517 4588 3523
rect 4740 3517 4892 3523
rect 5124 3517 5372 3523
rect 5428 3517 5484 3523
rect 5757 3523 5763 3537
rect 5956 3537 5964 3543
rect 5805 3524 5811 3536
rect 5572 3517 5772 3523
rect 5876 3517 5996 3523
rect 6004 3517 6044 3523
rect 2484 3497 2515 3503
rect 2525 3497 2540 3503
rect 1956 3477 2019 3483
rect 2036 3477 2099 3483
rect 148 3457 220 3463
rect 541 3463 547 3476
rect 541 3457 572 3463
rect 628 3457 652 3463
rect 724 3457 828 3463
rect 1028 3457 1100 3463
rect 1140 3457 1164 3463
rect 1188 3457 1356 3463
rect 1380 3457 1516 3463
rect 1540 3457 1724 3463
rect 1732 3457 1804 3463
rect 1812 3457 1964 3463
rect 2093 3463 2099 3477
rect 2116 3477 2172 3483
rect 2228 3477 2236 3483
rect 2260 3477 2428 3483
rect 2452 3477 2492 3483
rect 2509 3483 2515 3497
rect 2621 3497 2684 3503
rect 2509 3477 2572 3483
rect 2621 3483 2627 3497
rect 2845 3497 3340 3503
rect 2596 3477 2627 3483
rect 2845 3483 2851 3497
rect 3396 3497 3436 3503
rect 3460 3497 3628 3503
rect 3668 3497 3692 3503
rect 3700 3497 3708 3503
rect 3732 3497 3852 3503
rect 3940 3497 3948 3503
rect 3956 3497 4220 3503
rect 4228 3497 4556 3503
rect 4788 3497 4796 3503
rect 4804 3497 4844 3503
rect 4868 3497 4956 3503
rect 5476 3497 5532 3503
rect 5540 3497 5580 3503
rect 5588 3497 5628 3503
rect 5684 3497 5932 3503
rect 2644 3477 2851 3483
rect 2900 3477 2988 3483
rect 3357 3477 3459 3483
rect 3037 3464 3043 3476
rect 2093 3457 2204 3463
rect 2212 3457 2284 3463
rect 2292 3457 2316 3463
rect 2340 3457 2604 3463
rect 2621 3457 2700 3463
rect 180 3437 204 3443
rect 1796 3437 1836 3443
rect 1844 3437 1900 3443
rect 2068 3437 2092 3443
rect 2621 3443 2627 3457
rect 2756 3457 2876 3463
rect 3124 3457 3308 3463
rect 2429 3437 2627 3443
rect 932 3417 1004 3423
rect 1044 3417 1260 3423
rect 1332 3417 2124 3423
rect 2276 3417 2300 3423
rect 2429 3423 2435 3437
rect 2676 3437 2732 3443
rect 2749 3437 2972 3443
rect 2749 3423 2755 3437
rect 3060 3437 3132 3443
rect 3357 3443 3363 3477
rect 3453 3464 3459 3477
rect 3476 3477 3628 3483
rect 3636 3477 3660 3483
rect 3764 3477 4268 3483
rect 5092 3477 5132 3483
rect 5188 3477 5244 3483
rect 5268 3477 5484 3483
rect 5492 3477 5612 3483
rect 5620 3477 5644 3483
rect 5668 3477 5708 3483
rect 5732 3477 5852 3483
rect 5892 3477 5932 3483
rect 5972 3477 6076 3483
rect 3380 3457 3420 3463
rect 3556 3457 3564 3463
rect 3684 3457 3724 3463
rect 3764 3457 3788 3463
rect 3828 3457 3852 3463
rect 3860 3457 4588 3463
rect 4596 3457 4780 3463
rect 5284 3457 5340 3463
rect 5412 3457 5420 3463
rect 5428 3457 5724 3463
rect 5732 3457 5740 3463
rect 5748 3457 5964 3463
rect 5972 3457 6124 3463
rect 6132 3457 6156 3463
rect 3236 3437 3363 3443
rect 3380 3437 3468 3443
rect 3652 3437 3756 3443
rect 3780 3437 3916 3443
rect 3972 3437 4044 3443
rect 4132 3437 4172 3443
rect 4276 3437 4460 3443
rect 5284 3437 5420 3443
rect 5684 3437 5740 3443
rect 5748 3437 5964 3443
rect 5988 3437 6076 3443
rect 6100 3437 6124 3443
rect 6132 3437 6236 3443
rect 2324 3417 2435 3423
rect 2445 3417 2755 3423
rect 340 3397 492 3403
rect 548 3397 620 3403
rect 948 3397 956 3403
rect 1028 3397 1068 3403
rect 1124 3397 1180 3403
rect 1204 3397 1260 3403
rect 1332 3397 1436 3403
rect 1508 3397 1564 3403
rect 1652 3397 1708 3403
rect 1876 3397 1900 3403
rect 1972 3397 2076 3403
rect 2100 3397 2300 3403
rect 2356 3397 2380 3403
rect 2445 3403 2451 3417
rect 2836 3417 2908 3423
rect 2932 3417 2940 3423
rect 2996 3417 3084 3423
rect 3188 3417 3484 3423
rect 3636 3417 3660 3423
rect 3677 3417 3724 3423
rect 3112 3414 3160 3416
rect 3112 3406 3113 3414
rect 3122 3406 3123 3414
rect 3158 3406 3160 3414
rect 3112 3404 3160 3406
rect 3677 3404 3683 3417
rect 3748 3417 3980 3423
rect 4125 3417 4268 3423
rect 2420 3397 2451 3403
rect 2516 3397 2956 3403
rect 3188 3397 3235 3403
rect 1821 3384 1827 3396
rect 132 3377 364 3383
rect 372 3377 524 3383
rect 541 3377 684 3383
rect 196 3357 508 3363
rect 541 3363 547 3377
rect 884 3377 892 3383
rect 916 3377 940 3383
rect 1044 3377 1132 3383
rect 1236 3377 1244 3383
rect 1268 3377 1276 3383
rect 1428 3377 1820 3383
rect 1828 3377 2348 3383
rect 2356 3377 2364 3383
rect 2548 3377 2588 3383
rect 2628 3377 2636 3383
rect 2644 3377 2796 3383
rect 2852 3377 2924 3383
rect 2932 3377 2956 3383
rect 2980 3377 3148 3383
rect 3229 3383 3235 3397
rect 3252 3397 3420 3403
rect 3524 3397 3628 3403
rect 4125 3403 4131 3417
rect 5124 3417 5324 3423
rect 5844 3417 5916 3423
rect 6052 3417 6092 3423
rect 3700 3397 4131 3403
rect 4148 3397 4204 3403
rect 5236 3397 5292 3403
rect 5460 3397 5580 3403
rect 5748 3397 5772 3403
rect 5956 3397 5964 3403
rect 6004 3397 6060 3403
rect 3229 3377 3260 3383
rect 3284 3377 3292 3383
rect 3380 3377 3468 3383
rect 3508 3377 4300 3383
rect 4308 3377 4332 3383
rect 4340 3377 4748 3383
rect 4772 3377 4892 3383
rect 5364 3377 5436 3383
rect 5524 3377 5548 3383
rect 5828 3377 6012 3383
rect 6180 3377 6188 3383
rect 516 3357 547 3363
rect 564 3357 588 3363
rect 676 3357 828 3363
rect 852 3357 1068 3363
rect 1172 3357 1308 3363
rect 1332 3357 1532 3363
rect 1572 3357 1596 3363
rect 1716 3357 1852 3363
rect 1908 3357 1932 3363
rect 1988 3357 1996 3363
rect 2052 3357 2092 3363
rect 2116 3357 2156 3363
rect 2173 3357 2316 3363
rect 436 3337 556 3343
rect 596 3337 636 3343
rect 788 3337 908 3343
rect 916 3337 1004 3343
rect 1044 3337 1244 3343
rect 2173 3343 2179 3357
rect 2372 3357 2572 3363
rect 1540 3337 2179 3343
rect 2212 3337 2252 3343
rect 2260 3337 2355 3343
rect 2349 3324 2355 3337
rect 2388 3337 2412 3343
rect 2477 3343 2483 3357
rect 2509 3343 2515 3357
rect 2612 3357 2668 3363
rect 2788 3357 2876 3363
rect 2996 3357 3084 3363
rect 3252 3357 3372 3363
rect 3460 3357 3532 3363
rect 3556 3357 3580 3363
rect 3620 3357 3660 3363
rect 3700 3357 3756 3363
rect 3780 3357 3804 3363
rect 3828 3357 5244 3363
rect 5252 3357 5292 3363
rect 5396 3357 5452 3363
rect 5460 3357 5548 3363
rect 5604 3357 5628 3363
rect 5652 3357 5708 3363
rect 5748 3357 6124 3363
rect 6132 3357 6140 3363
rect 2573 3344 2579 3356
rect 2477 3337 2572 3343
rect 2612 3337 2636 3343
rect 2653 3337 2828 3343
rect 180 3317 227 3323
rect 221 3264 227 3317
rect 276 3317 300 3323
rect 484 3317 604 3323
rect 612 3317 620 3323
rect 644 3317 684 3323
rect 724 3317 764 3323
rect 772 3317 828 3323
rect 852 3317 899 3323
rect 500 3297 588 3303
rect 676 3297 716 3303
rect 756 3297 844 3303
rect 468 3277 556 3283
rect 564 3277 588 3283
rect 893 3283 899 3317
rect 916 3317 972 3323
rect 996 3317 1052 3323
rect 1092 3317 1116 3323
rect 1172 3317 1276 3323
rect 1428 3317 1500 3323
rect 1588 3317 1676 3323
rect 1716 3317 1756 3323
rect 1764 3317 1804 3323
rect 1844 3317 1884 3323
rect 1892 3317 2124 3323
rect 2132 3317 2188 3323
rect 2212 3317 2252 3323
rect 2276 3317 2316 3323
rect 2356 3317 2412 3323
rect 2436 3317 2524 3323
rect 2653 3323 2659 3337
rect 2884 3337 2956 3343
rect 3188 3337 3212 3343
rect 3428 3337 3468 3343
rect 3508 3337 3532 3343
rect 3556 3337 3820 3343
rect 3892 3337 4060 3343
rect 4084 3337 4108 3343
rect 4116 3337 4156 3343
rect 4244 3337 4348 3343
rect 4484 3337 4604 3343
rect 4612 3337 4732 3343
rect 4740 3337 4956 3343
rect 5172 3337 5180 3343
rect 5236 3337 5644 3343
rect 5748 3337 5820 3343
rect 5844 3337 5884 3343
rect 5908 3337 5964 3343
rect 6013 3337 6028 3343
rect 6013 3324 6019 3337
rect 6068 3337 6188 3343
rect 2548 3317 2659 3323
rect 2676 3317 2748 3323
rect 2948 3317 3084 3323
rect 3172 3317 3276 3323
rect 3348 3317 3372 3323
rect 3428 3317 3500 3323
rect 3636 3317 3644 3323
rect 3652 3317 3692 3323
rect 3860 3317 3884 3323
rect 3924 3317 4172 3323
rect 4276 3317 4316 3323
rect 4324 3317 4492 3323
rect 4500 3317 4780 3323
rect 4804 3317 4844 3323
rect 4868 3317 5004 3323
rect 5060 3317 5116 3323
rect 5172 3317 5324 3323
rect 5348 3317 5420 3323
rect 5437 3317 5516 3323
rect 980 3297 1164 3303
rect 1172 3297 1180 3303
rect 1188 3297 1292 3303
rect 1364 3297 1388 3303
rect 1460 3297 1676 3303
rect 1940 3297 1964 3303
rect 2052 3297 2060 3303
rect 2164 3297 2444 3303
rect 2500 3297 2604 3303
rect 2644 3297 2668 3303
rect 2724 3297 2988 3303
rect 3012 3297 3052 3303
rect 3092 3297 3100 3303
rect 3108 3297 3180 3303
rect 3188 3297 3212 3303
rect 3252 3297 3356 3303
rect 3380 3297 3820 3303
rect 4036 3297 4268 3303
rect 4324 3297 4412 3303
rect 4436 3297 4844 3303
rect 4900 3297 5084 3303
rect 5124 3297 5164 3303
rect 5204 3297 5244 3303
rect 5332 3297 5340 3303
rect 5437 3303 5443 3317
rect 5540 3317 5596 3323
rect 5620 3317 5900 3323
rect 6036 3317 6252 3323
rect 5364 3297 5443 3303
rect 5508 3297 5580 3303
rect 5588 3297 5660 3303
rect 5812 3297 5900 3303
rect 5940 3297 5980 3303
rect 5988 3297 6076 3303
rect 6084 3297 6140 3303
rect 6164 3297 6188 3303
rect 6196 3297 6220 3303
rect 893 3277 1068 3283
rect 1108 3277 1404 3283
rect 1412 3277 1548 3283
rect 1556 3277 2108 3283
rect 2116 3277 3932 3283
rect 3940 3277 4636 3283
rect 5268 3277 5436 3283
rect 5476 3277 5948 3283
rect 6116 3277 6124 3283
rect 6212 3277 6252 3283
rect 532 3257 812 3263
rect 884 3257 1356 3263
rect 1396 3257 1420 3263
rect 1444 3257 1548 3263
rect 1668 3257 1708 3263
rect 1732 3257 1740 3263
rect 1780 3257 1820 3263
rect 1908 3257 1932 3263
rect 1972 3257 2028 3263
rect 2068 3257 2140 3263
rect 2164 3257 2284 3263
rect 2340 3257 2348 3263
rect 2372 3257 2508 3263
rect 2532 3257 2588 3263
rect 2612 3257 2700 3263
rect 2740 3257 2828 3263
rect 2852 3257 2860 3263
rect 2932 3257 3212 3263
rect 3220 3257 3228 3263
rect 3325 3257 3420 3263
rect 20 3237 467 3243
rect 276 3217 348 3223
rect 436 3217 444 3223
rect 461 3223 467 3237
rect 612 3237 684 3243
rect 724 3237 876 3243
rect 1012 3237 1068 3243
rect 1092 3237 1132 3243
rect 1149 3237 1900 3243
rect 1149 3223 1155 3237
rect 1924 3237 2092 3243
rect 2132 3237 2796 3243
rect 2836 3237 2876 3243
rect 2884 3237 3004 3243
rect 3325 3243 3331 3257
rect 3476 3257 4476 3263
rect 5364 3257 5388 3263
rect 5876 3257 6028 3263
rect 6052 3257 6108 3263
rect 3092 3237 3331 3243
rect 3364 3237 3388 3243
rect 3444 3237 3756 3243
rect 3780 3237 3804 3243
rect 3860 3237 3964 3243
rect 4100 3237 5100 3243
rect 5396 3237 5580 3243
rect 5956 3237 6188 3243
rect 461 3217 1155 3223
rect 1364 3217 1516 3223
rect 1700 3217 1724 3223
rect 1732 3217 1772 3223
rect 1796 3217 1932 3223
rect 2148 3217 2204 3223
rect 2292 3217 2460 3223
rect 2500 3217 2508 3223
rect 2557 3217 2700 3223
rect 1576 3214 1624 3216
rect 1576 3206 1577 3214
rect 1586 3206 1587 3214
rect 1622 3206 1624 3214
rect 1576 3204 1624 3206
rect 148 3197 412 3203
rect 548 3197 588 3203
rect 596 3197 844 3203
rect 884 3197 1116 3203
rect 1236 3197 1244 3203
rect 1268 3197 1420 3203
rect 1476 3197 1516 3203
rect 1668 3197 2012 3203
rect 2020 3197 2220 3203
rect 2557 3203 2563 3217
rect 2788 3217 2812 3223
rect 2868 3217 2892 3223
rect 2916 3217 2940 3223
rect 2980 3217 3372 3223
rect 3412 3217 4108 3223
rect 4664 3214 4712 3216
rect 4664 3206 4665 3214
rect 4674 3206 4675 3214
rect 4710 3206 4712 3214
rect 4664 3204 4712 3206
rect 2228 3197 2563 3203
rect 2580 3197 2604 3203
rect 2612 3197 3548 3203
rect 3748 3197 3852 3203
rect 3876 3197 3980 3203
rect 4020 3197 4124 3203
rect 4148 3197 4508 3203
rect 5396 3197 5404 3203
rect 196 3177 588 3183
rect 852 3177 1036 3183
rect 1156 3177 1292 3183
rect 1316 3177 1475 3183
rect 148 3157 204 3163
rect 372 3157 412 3163
rect 420 3157 579 3163
rect 324 3137 428 3143
rect 436 3137 460 3143
rect 573 3143 579 3157
rect 596 3157 604 3163
rect 740 3157 780 3163
rect 948 3157 1196 3163
rect 1204 3157 1212 3163
rect 1236 3157 1324 3163
rect 1469 3163 1475 3177
rect 1492 3177 1692 3183
rect 1716 3177 1900 3183
rect 2100 3177 2380 3183
rect 2404 3177 2732 3183
rect 2804 3177 3036 3183
rect 3108 3177 3244 3183
rect 3268 3177 3436 3183
rect 3476 3177 3484 3183
rect 3508 3177 4332 3183
rect 5204 3177 5804 3183
rect 5812 3177 5948 3183
rect 6052 3177 6092 3183
rect 1469 3157 2156 3163
rect 2292 3157 2316 3163
rect 2333 3157 2428 3163
rect 573 3137 716 3143
rect 1012 3137 1244 3143
rect 1300 3137 1523 3143
rect 557 3124 563 3136
rect 100 3117 220 3123
rect 356 3117 460 3123
rect 468 3117 492 3123
rect 580 3117 588 3123
rect 660 3117 716 3123
rect 724 3117 908 3123
rect 948 3117 988 3123
rect 996 3117 1068 3123
rect 1156 3117 1171 3123
rect 1165 3104 1171 3117
rect 1204 3117 1228 3123
rect 1252 3117 1260 3123
rect 1428 3117 1500 3123
rect 1517 3123 1523 3137
rect 1540 3137 1580 3143
rect 1652 3137 1788 3143
rect 1828 3137 1843 3143
rect 1517 3117 1548 3123
rect 1572 3117 1644 3123
rect 1684 3117 1708 3123
rect 1837 3123 1843 3137
rect 1876 3137 1900 3143
rect 1940 3137 1964 3143
rect 2004 3137 2028 3143
rect 2333 3143 2339 3157
rect 2516 3157 2636 3163
rect 2660 3157 2668 3163
rect 2740 3157 2972 3163
rect 3396 3157 3404 3163
rect 3428 3157 3660 3163
rect 3684 3157 3692 3163
rect 3828 3157 4092 3163
rect 4148 3157 5084 3163
rect 5092 3157 5164 3163
rect 5332 3157 5756 3163
rect 5908 3157 5932 3163
rect 5972 3157 5996 3163
rect 6036 3157 6092 3163
rect 2068 3137 2339 3143
rect 2436 3137 2508 3143
rect 2548 3137 2748 3143
rect 2868 3137 2940 3143
rect 2964 3137 3052 3143
rect 3156 3137 3196 3143
rect 3348 3137 3772 3143
rect 3796 3137 3820 3143
rect 3860 3137 3980 3143
rect 4004 3137 4028 3143
rect 4052 3137 4172 3143
rect 4676 3137 4796 3143
rect 5508 3137 5548 3143
rect 5604 3137 5628 3143
rect 5924 3137 5980 3143
rect 6164 3137 6220 3143
rect 1837 3117 1868 3123
rect 1892 3117 1980 3123
rect 1997 3117 2060 3123
rect 228 3097 236 3103
rect 260 3097 284 3103
rect 340 3097 524 3103
rect 580 3097 620 3103
rect 820 3097 908 3103
rect 980 3097 988 3103
rect 1028 3097 1036 3103
rect 580 3077 588 3083
rect 596 3077 620 3083
rect 692 3077 748 3083
rect 868 3077 876 3083
rect 916 3077 1020 3083
rect 1181 3083 1187 3116
rect 1204 3097 1244 3103
rect 1268 3097 1276 3103
rect 1396 3097 1484 3103
rect 1524 3097 1564 3103
rect 1604 3097 1740 3103
rect 1780 3097 1836 3103
rect 1997 3103 2003 3117
rect 2132 3117 2259 3123
rect 1972 3097 2003 3103
rect 2068 3097 2124 3103
rect 2164 3097 2204 3103
rect 2253 3103 2259 3117
rect 2276 3117 2364 3123
rect 2388 3117 2444 3123
rect 2461 3117 2540 3123
rect 2461 3103 2467 3117
rect 2596 3117 2860 3123
rect 2980 3117 3084 3123
rect 3380 3117 3420 3123
rect 3460 3117 3484 3123
rect 3620 3117 3708 3123
rect 3732 3117 3884 3123
rect 3924 3117 4108 3123
rect 4132 3117 4156 3123
rect 4180 3117 4188 3123
rect 4788 3117 4844 3123
rect 5188 3117 5276 3123
rect 5316 3117 5420 3123
rect 5540 3117 5596 3123
rect 5812 3117 5884 3123
rect 5908 3117 6060 3123
rect 6068 3117 6124 3123
rect 6164 3117 6188 3123
rect 6196 3117 6236 3123
rect 2253 3097 2467 3103
rect 2484 3097 2636 3103
rect 2788 3097 2796 3103
rect 2836 3097 3075 3103
rect 1156 3077 1187 3083
rect 1220 3077 1388 3083
rect 1453 3077 1532 3083
rect 205 3064 211 3076
rect 564 3057 700 3063
rect 772 3057 780 3063
rect 884 3057 924 3063
rect 932 3057 956 3063
rect 980 3057 1308 3063
rect 1453 3063 1459 3077
rect 1556 3077 1660 3083
rect 1748 3077 1756 3083
rect 1812 3077 1884 3083
rect 1940 3077 2268 3083
rect 2356 3077 2380 3083
rect 2404 3077 2460 3083
rect 2516 3077 2572 3083
rect 2612 3077 2620 3083
rect 2644 3077 2684 3083
rect 2701 3077 2732 3083
rect 1332 3057 1459 3063
rect 1476 3057 1500 3063
rect 1508 3057 1532 3063
rect 1620 3057 1635 3063
rect 292 3037 300 3043
rect 308 3037 636 3043
rect 1140 3037 1180 3043
rect 500 3017 508 3023
rect 628 3017 844 3023
rect 884 3017 924 3023
rect 948 3017 972 3023
rect 1012 3017 1084 3023
rect 1124 3017 1388 3023
rect 1444 3017 1580 3023
rect 1629 3023 1635 3057
rect 1652 3057 1692 3063
rect 1700 3057 1708 3063
rect 1748 3057 1788 3063
rect 1844 3057 1852 3063
rect 1908 3057 1964 3063
rect 2004 3057 2028 3063
rect 2052 3057 2076 3063
rect 2100 3057 2172 3063
rect 2260 3057 2284 3063
rect 2356 3057 2364 3063
rect 2701 3063 2707 3077
rect 2804 3077 2860 3083
rect 2996 3077 3020 3083
rect 3069 3083 3075 3097
rect 3092 3097 3532 3103
rect 3613 3097 3948 3103
rect 3069 3077 3100 3083
rect 3188 3077 3228 3083
rect 3236 3077 3276 3083
rect 3348 3077 3532 3083
rect 3613 3083 3619 3097
rect 4052 3097 4300 3103
rect 4356 3097 4428 3103
rect 4532 3097 4876 3103
rect 5012 3097 5052 3103
rect 5220 3097 5276 3103
rect 5428 3097 5452 3103
rect 5556 3097 5644 3103
rect 5716 3097 5836 3103
rect 5844 3097 5916 3103
rect 5940 3097 5980 3103
rect 6164 3097 6188 3103
rect 6212 3097 6284 3103
rect 3588 3077 3619 3083
rect 3668 3077 3692 3083
rect 3716 3077 3772 3083
rect 3796 3077 3868 3083
rect 3892 3077 3932 3083
rect 3965 3077 4060 3083
rect 2452 3057 2707 3063
rect 2740 3057 2876 3063
rect 3357 3057 3388 3063
rect 1668 3037 1708 3043
rect 1716 3037 1820 3043
rect 1844 3037 2028 3043
rect 2052 3037 2156 3043
rect 2260 3037 2396 3043
rect 2420 3037 2444 3043
rect 2580 3037 2620 3043
rect 2676 3037 2796 3043
rect 2813 3037 2972 3043
rect 1629 3017 1676 3023
rect 1764 3017 1900 3023
rect 1940 3017 1980 3023
rect 2004 3017 2188 3023
rect 2244 3017 2268 3023
rect 2292 3017 2300 3023
rect 2516 3017 2588 3023
rect 2612 3017 2652 3023
rect 2813 3023 2819 3037
rect 2996 3037 3020 3043
rect 3076 3037 3164 3043
rect 3181 3043 3187 3056
rect 3181 3037 3203 3043
rect 2804 3017 2819 3023
rect 2916 3017 2940 3023
rect 3197 3023 3203 3037
rect 3220 3037 3244 3043
rect 3357 3043 3363 3057
rect 3412 3057 3436 3063
rect 3453 3057 3596 3063
rect 3252 3037 3363 3043
rect 3453 3043 3459 3057
rect 3965 3063 3971 3077
rect 4084 3077 4220 3083
rect 4228 3077 4268 3083
rect 4308 3077 4332 3083
rect 4420 3077 4460 3083
rect 4708 3077 4732 3083
rect 5172 3077 5324 3083
rect 5428 3077 5452 3083
rect 5476 3077 5516 3083
rect 5524 3077 5676 3083
rect 5780 3077 5884 3083
rect 5908 3077 5932 3083
rect 5940 3077 6220 3083
rect 3652 3057 3971 3063
rect 3988 3057 5187 3063
rect 3380 3037 3459 3043
rect 3476 3037 3500 3043
rect 3588 3037 3836 3043
rect 3876 3037 4204 3043
rect 4404 3037 4428 3043
rect 4468 3037 4508 3043
rect 4532 3037 4732 3043
rect 5181 3043 5187 3057
rect 5332 3057 5340 3063
rect 5412 3057 5420 3063
rect 5428 3057 5436 3063
rect 5492 3057 5635 3063
rect 5181 3037 5532 3043
rect 5629 3043 5635 3057
rect 5652 3057 5676 3063
rect 5684 3057 5980 3063
rect 6052 3057 6076 3063
rect 6116 3057 6140 3063
rect 6148 3057 6156 3063
rect 5629 3037 5724 3043
rect 5844 3037 6044 3043
rect 6148 3037 6236 3043
rect 3197 3017 3228 3023
rect 3316 3017 3340 3023
rect 3364 3017 4140 3023
rect 4212 3017 4284 3023
rect 4356 3017 4428 3023
rect 4500 3017 5292 3023
rect 5300 3017 5388 3023
rect 5556 3017 5788 3023
rect 6132 3017 6172 3023
rect 3112 3014 3160 3016
rect 3112 3006 3113 3014
rect 3122 3006 3123 3014
rect 3158 3006 3160 3014
rect 3112 3004 3160 3006
rect 548 2997 588 3003
rect 724 2997 1452 3003
rect 1524 2997 1644 3003
rect 1908 2997 2044 3003
rect 2084 2997 2140 3003
rect 2164 2997 2188 3003
rect 2212 2997 2348 3003
rect 2372 2997 2524 3003
rect 2548 2997 2556 3003
rect 2612 2997 2732 3003
rect 2756 2997 2812 3003
rect 2868 2997 2892 3003
rect 2932 2997 2956 3003
rect 2996 2997 3004 3003
rect 3268 2997 3340 3003
rect 3348 2997 3404 3003
rect 3444 2997 3660 3003
rect 3764 2997 4012 3003
rect 4084 2997 5228 3003
rect 5268 2997 5667 3003
rect 244 2977 348 2983
rect 692 2977 1212 2983
rect 1236 2977 1420 2983
rect 1460 2977 3452 2983
rect 3460 2977 3852 2983
rect 3908 2977 3932 2983
rect 4100 2977 4284 2983
rect 4292 2977 4652 2983
rect 5661 2983 5667 2997
rect 5684 2997 5868 3003
rect 6180 2997 6268 3003
rect 5661 2977 5692 2983
rect 6260 2977 6275 2983
rect 36 2957 332 2963
rect 548 2957 604 2963
rect 660 2957 700 2963
rect 708 2957 732 2963
rect 788 2957 796 2963
rect 820 2957 1052 2963
rect 1060 2957 1148 2963
rect 1172 2957 1388 2963
rect 1405 2957 1612 2963
rect 340 2937 380 2943
rect 516 2937 556 2943
rect 884 2937 1004 2943
rect 1076 2937 1116 2943
rect 1220 2937 1308 2943
rect 1316 2937 1324 2943
rect 1405 2943 1411 2957
rect 1684 2957 1724 2963
rect 1812 2957 1932 2963
rect 1940 2957 1996 2963
rect 2036 2957 2188 2963
rect 2212 2957 2252 2963
rect 2260 2957 2300 2963
rect 2324 2957 2476 2963
rect 2484 2957 2668 2963
rect 2740 2957 2764 2963
rect 2788 2957 2796 2963
rect 2932 2957 3059 2963
rect 1380 2937 1411 2943
rect 1428 2937 2188 2943
rect 2228 2937 2268 2943
rect 2356 2937 2444 2943
rect 2580 2937 2636 2943
rect 2772 2937 2892 2943
rect 2980 2937 3036 2943
rect 3053 2943 3059 2957
rect 3076 2957 3084 2963
rect 3124 2957 3180 2963
rect 3204 2957 3308 2963
rect 3316 2957 3356 2963
rect 3396 2957 3404 2963
rect 3604 2957 3635 2963
rect 3053 2937 3260 2943
rect 3284 2937 3308 2943
rect 3332 2937 3372 2943
rect 3444 2937 3612 2943
rect 3629 2943 3635 2957
rect 3684 2957 3724 2963
rect 3732 2957 4044 2963
rect 3629 2937 3692 2943
rect 3732 2937 3964 2943
rect 4077 2943 4083 2976
rect 6269 2964 6275 2977
rect 4372 2957 4380 2963
rect 4580 2957 4652 2963
rect 4660 2957 4972 2963
rect 5220 2957 5228 2963
rect 5348 2957 5372 2963
rect 5444 2957 5484 2963
rect 5524 2957 5548 2963
rect 5572 2957 5644 2963
rect 5684 2957 5740 2963
rect 5988 2957 6076 2963
rect 6196 2957 6252 2963
rect 4068 2937 4083 2943
rect 4180 2937 4236 2943
rect 4276 2937 4316 2943
rect 4324 2937 4540 2943
rect 4644 2937 4684 2943
rect 4740 2937 4908 2943
rect 4916 2937 5036 2943
rect 5156 2937 5292 2943
rect 5428 2937 5644 2943
rect 5652 2937 5692 2943
rect 5812 2937 6028 2943
rect 6068 2937 6076 2943
rect 6084 2937 6124 2943
rect 6132 2937 6220 2943
rect 1037 2924 1043 2936
rect 5741 2924 5747 2936
rect 68 2917 156 2923
rect 548 2917 572 2923
rect 580 2917 748 2923
rect 852 2917 1020 2923
rect 1092 2917 1132 2923
rect 1140 2917 1187 2923
rect 397 2904 403 2916
rect 20 2897 156 2903
rect 164 2897 220 2903
rect 372 2897 396 2903
rect 420 2897 732 2903
rect 884 2897 908 2903
rect 964 2897 988 2903
rect 1044 2897 1100 2903
rect 1140 2897 1164 2903
rect 1181 2903 1187 2917
rect 1252 2917 1260 2923
rect 1469 2917 1532 2923
rect 1181 2897 1340 2903
rect 1469 2903 1475 2917
rect 1540 2917 1587 2923
rect 1421 2897 1475 2903
rect 292 2877 460 2883
rect 477 2877 716 2883
rect 84 2857 140 2863
rect 148 2857 188 2863
rect 196 2857 252 2863
rect 477 2863 483 2877
rect 724 2877 956 2883
rect 1076 2877 1180 2883
rect 1421 2883 1427 2897
rect 1508 2897 1532 2903
rect 1556 2897 1564 2903
rect 1581 2903 1587 2917
rect 1604 2917 1740 2923
rect 1828 2917 1868 2923
rect 1876 2917 1900 2923
rect 2452 2917 2508 2923
rect 2525 2917 2732 2923
rect 1581 2897 1756 2903
rect 1844 2897 2092 2903
rect 2125 2897 2156 2903
rect 1188 2877 1427 2883
rect 1444 2877 1772 2883
rect 1860 2877 1868 2883
rect 1892 2877 1932 2883
rect 2004 2877 2092 2883
rect 2125 2883 2131 2897
rect 2180 2897 2284 2903
rect 2340 2897 2364 2903
rect 2388 2897 2435 2903
rect 2116 2877 2131 2883
rect 2196 2877 2220 2883
rect 2429 2883 2435 2897
rect 2525 2903 2531 2917
rect 2756 2917 2851 2923
rect 2516 2897 2531 2903
rect 2548 2897 2620 2903
rect 2676 2897 2684 2903
rect 2845 2903 2851 2917
rect 2916 2917 2940 2923
rect 2996 2917 3020 2923
rect 3060 2917 3100 2923
rect 3236 2917 3276 2923
rect 3284 2917 3420 2923
rect 3444 2917 3500 2923
rect 3508 2917 3724 2923
rect 3796 2917 3916 2923
rect 3956 2917 3980 2923
rect 4020 2917 4092 2923
rect 4132 2917 4348 2923
rect 4372 2917 4396 2923
rect 4532 2917 4588 2923
rect 4596 2917 4636 2923
rect 4868 2917 5020 2923
rect 5076 2917 5260 2923
rect 5284 2917 5612 2923
rect 5620 2917 5628 2923
rect 5645 2917 5740 2923
rect 2692 2897 2787 2903
rect 2845 2897 3244 2903
rect 2429 2877 2460 2883
rect 2564 2877 2764 2883
rect 2781 2883 2787 2897
rect 3284 2897 3532 2903
rect 3556 2897 3596 2903
rect 3620 2897 3644 2903
rect 3668 2897 3708 2903
rect 3716 2897 3916 2903
rect 3924 2897 3948 2903
rect 4020 2897 4300 2903
rect 5124 2897 5164 2903
rect 5172 2897 5196 2903
rect 5645 2903 5651 2917
rect 6148 2917 6172 2923
rect 6212 2917 6236 2923
rect 5220 2897 5651 2903
rect 5700 2897 5788 2903
rect 5972 2897 5996 2903
rect 6148 2897 6188 2903
rect 2781 2877 2988 2883
rect 3044 2877 3052 2883
rect 3076 2877 3180 2883
rect 3204 2877 3340 2883
rect 3668 2877 4012 2883
rect 4020 2877 4892 2883
rect 5028 2877 5116 2883
rect 5476 2877 5516 2883
rect 5812 2877 5820 2883
rect 6020 2877 6108 2883
rect 404 2857 483 2863
rect 596 2857 908 2863
rect 980 2857 1132 2863
rect 1428 2857 1612 2863
rect 1636 2857 1660 2863
rect 1684 2857 1708 2863
rect 1748 2857 1804 2863
rect 1844 2857 2140 2863
rect 2164 2857 2252 2863
rect 2340 2857 2508 2863
rect 2548 2857 2636 2863
rect 2900 2857 2988 2863
rect 3028 2857 3052 2863
rect 3069 2857 3116 2863
rect 324 2837 524 2843
rect 532 2837 604 2843
rect 612 2837 1100 2843
rect 1172 2837 1228 2843
rect 1300 2837 1772 2843
rect 1876 2837 1996 2843
rect 2020 2837 2044 2843
rect 2116 2837 2284 2843
rect 2292 2837 2508 2843
rect 2708 2837 2796 2843
rect 2884 2837 2892 2843
rect 3069 2843 3075 2857
rect 3140 2857 3372 2863
rect 3476 2857 3548 2863
rect 3604 2857 3804 2863
rect 3812 2857 3868 2863
rect 4068 2857 4140 2863
rect 5236 2857 5276 2863
rect 5284 2857 5324 2863
rect 5508 2857 5580 2863
rect 5588 2857 5724 2863
rect 5892 2857 5996 2863
rect 6004 2857 6028 2863
rect 2996 2837 3075 2843
rect 3092 2837 3116 2843
rect 3236 2837 3244 2843
rect 3268 2837 3324 2843
rect 3364 2837 3388 2843
rect 3444 2837 3452 2843
rect 3565 2837 3612 2843
rect 244 2817 652 2823
rect 660 2817 844 2823
rect 900 2817 924 2823
rect 964 2817 1116 2823
rect 1156 2817 1180 2823
rect 1268 2817 1548 2823
rect 1684 2817 1788 2823
rect 1812 2817 1948 2823
rect 1972 2817 2124 2823
rect 2164 2817 2204 2823
rect 2292 2817 2428 2823
rect 2452 2817 2588 2823
rect 2756 2817 2860 2823
rect 3044 2817 3164 2823
rect 3565 2823 3571 2837
rect 3668 2837 4620 2843
rect 4644 2837 4684 2843
rect 5508 2837 5708 2843
rect 5780 2837 6236 2843
rect 3252 2817 3571 2823
rect 3588 2817 4620 2823
rect 5684 2817 5804 2823
rect 5876 2817 6252 2823
rect 1576 2814 1624 2816
rect 1576 2806 1577 2814
rect 1586 2806 1587 2814
rect 1622 2806 1624 2814
rect 1576 2804 1624 2806
rect 4664 2814 4712 2816
rect 4664 2806 4665 2814
rect 4674 2806 4675 2814
rect 4710 2806 4712 2814
rect 4664 2804 4712 2806
rect 500 2797 572 2803
rect 916 2797 972 2803
rect 1076 2797 1228 2803
rect 1332 2797 1356 2803
rect 1373 2797 1452 2803
rect 132 2777 140 2783
rect 148 2777 220 2783
rect 228 2777 668 2783
rect 900 2777 1196 2783
rect 1204 2777 1260 2783
rect 1373 2783 1379 2797
rect 1492 2797 1516 2803
rect 1700 2797 1804 2803
rect 2164 2797 3052 2803
rect 3188 2797 3516 2803
rect 3572 2797 3772 2803
rect 3796 2797 3836 2803
rect 3860 2797 3884 2803
rect 3892 2797 3900 2803
rect 3924 2797 3948 2803
rect 4020 2797 4076 2803
rect 4164 2797 4300 2803
rect 5604 2797 5628 2803
rect 5636 2797 6012 2803
rect 6164 2797 6188 2803
rect 1316 2777 1379 2783
rect 1396 2777 1452 2783
rect 1524 2777 1756 2783
rect 1780 2777 2179 2783
rect 180 2757 220 2763
rect 244 2757 412 2763
rect 532 2757 556 2763
rect 676 2757 892 2763
rect 948 2757 1212 2763
rect 1236 2757 1324 2763
rect 1460 2757 1532 2763
rect 1540 2757 1676 2763
rect 1716 2757 1788 2763
rect 1812 2757 2156 2763
rect 2173 2763 2179 2777
rect 2196 2777 2444 2783
rect 2484 2777 2540 2783
rect 2573 2777 2716 2783
rect 2173 2757 2348 2763
rect 2388 2757 2492 2763
rect 2573 2744 2579 2777
rect 2740 2777 3068 2783
rect 3108 2777 3164 2783
rect 3220 2777 3292 2783
rect 3316 2777 3532 2783
rect 3732 2777 3756 2783
rect 3780 2777 4044 2783
rect 4244 2777 4284 2783
rect 4628 2777 5276 2783
rect 5332 2777 5468 2783
rect 5684 2777 5852 2783
rect 5860 2777 6156 2783
rect 2660 2757 2684 2763
rect 2708 2757 2755 2763
rect 100 2737 252 2743
rect 372 2737 428 2743
rect 452 2737 556 2743
rect 564 2737 940 2743
rect 964 2737 1091 2743
rect 164 2717 188 2723
rect 340 2717 540 2723
rect 596 2717 636 2723
rect 708 2717 748 2723
rect 884 2717 908 2723
rect 916 2717 956 2723
rect 1085 2704 1091 2737
rect 1124 2737 1148 2743
rect 1188 2737 1260 2743
rect 1524 2737 1548 2743
rect 1572 2737 1644 2743
rect 1661 2737 1740 2743
rect 1108 2717 1164 2723
rect 1172 2717 1228 2723
rect 1661 2723 1667 2737
rect 1780 2737 1820 2743
rect 1837 2737 1964 2743
rect 1396 2717 1667 2723
rect 1837 2723 1843 2737
rect 2004 2737 2220 2743
rect 2260 2737 2556 2743
rect 2596 2737 2732 2743
rect 2749 2743 2755 2757
rect 2820 2757 2924 2763
rect 2948 2757 3004 2763
rect 3028 2760 3356 2763
rect 3021 2757 3356 2760
rect 3380 2757 3564 2763
rect 3604 2757 3740 2763
rect 3764 2757 3948 2763
rect 3965 2757 4076 2763
rect 2749 2737 2764 2743
rect 2804 2737 3004 2743
rect 3021 2740 3052 2743
rect 3028 2737 3052 2740
rect 3076 2737 3187 2743
rect 1828 2717 1843 2723
rect 2132 2717 2188 2723
rect 2372 2717 2604 2723
rect 2660 2717 2764 2723
rect 2852 2717 2860 2723
rect 2900 2717 2924 2723
rect 2948 2717 2972 2723
rect 3028 2717 3084 2723
rect 3101 2717 3148 2723
rect 1677 2704 1683 2716
rect 84 2697 172 2703
rect 276 2697 364 2703
rect 420 2697 428 2703
rect 468 2697 620 2703
rect 628 2697 956 2703
rect 1021 2697 1052 2703
rect 180 2677 220 2683
rect 372 2677 380 2683
rect 500 2677 508 2683
rect 532 2677 716 2683
rect 1021 2683 1027 2697
rect 1108 2697 1564 2703
rect 1757 2703 1763 2716
rect 1684 2697 1731 2703
rect 1757 2697 1836 2703
rect 868 2677 1027 2683
rect 1044 2677 1052 2683
rect 1172 2677 1244 2683
rect 1268 2677 1292 2683
rect 1300 2677 1388 2683
rect 1428 2677 1468 2683
rect 1492 2677 1548 2683
rect 1556 2677 1692 2683
rect 1725 2683 1731 2697
rect 1860 2697 1884 2703
rect 1917 2703 1923 2716
rect 1917 2697 1996 2703
rect 2084 2697 2220 2703
rect 2228 2697 2444 2703
rect 2500 2697 2524 2703
rect 2548 2697 2684 2703
rect 2708 2697 2748 2703
rect 2772 2697 2908 2703
rect 3101 2703 3107 2717
rect 3181 2723 3187 2737
rect 3204 2737 3260 2743
rect 3268 2737 3276 2743
rect 3300 2737 3308 2743
rect 3444 2737 3788 2743
rect 3965 2743 3971 2757
rect 4292 2757 4524 2763
rect 4628 2757 5724 2763
rect 5748 2757 5804 2763
rect 5892 2757 5932 2763
rect 3828 2737 3971 2743
rect 3988 2737 4044 2743
rect 4084 2737 4396 2743
rect 4500 2737 5500 2743
rect 5524 2737 5580 2743
rect 5748 2737 5772 2743
rect 5908 2737 5980 2743
rect 6132 2737 6140 2743
rect 3181 2717 3228 2723
rect 3236 2717 3244 2723
rect 3300 2717 3404 2723
rect 3460 2717 3516 2723
rect 3556 2717 3596 2723
rect 3604 2717 3852 2723
rect 3860 2717 4796 2723
rect 5156 2717 5340 2723
rect 5572 2717 5580 2723
rect 5620 2717 5628 2723
rect 5716 2717 5868 2723
rect 5885 2717 5932 2723
rect 2996 2697 3107 2703
rect 3124 2697 3596 2703
rect 3636 2697 3683 2703
rect 1725 2677 1756 2683
rect 1780 2677 1852 2683
rect 1924 2677 1948 2683
rect 1956 2677 1964 2683
rect 2004 2677 2188 2683
rect 2212 2677 2300 2683
rect 2308 2677 2316 2683
rect 2452 2677 2476 2683
rect 2516 2677 2652 2683
rect 2692 2677 2748 2683
rect 2829 2677 2956 2683
rect 468 2657 572 2663
rect 724 2657 1187 2663
rect 436 2637 492 2643
rect 500 2637 1164 2643
rect 1181 2643 1187 2657
rect 1204 2657 1228 2663
rect 1252 2657 1276 2663
rect 1300 2657 1372 2663
rect 1428 2657 1484 2663
rect 1508 2657 1596 2663
rect 1700 2657 1795 2663
rect 1181 2637 1276 2643
rect 1380 2637 1404 2643
rect 1476 2637 1484 2643
rect 1508 2637 1596 2643
rect 1620 2637 1708 2643
rect 1732 2637 1772 2643
rect 1789 2643 1795 2657
rect 1812 2657 1868 2663
rect 1908 2657 2044 2663
rect 2100 2657 2188 2663
rect 2260 2657 2275 2663
rect 1789 2637 1804 2643
rect 1828 2637 1836 2643
rect 1892 2637 1964 2643
rect 2036 2637 2236 2643
rect 2269 2643 2275 2657
rect 2356 2657 2428 2663
rect 2468 2657 2556 2663
rect 2612 2657 2636 2663
rect 2676 2657 2684 2663
rect 2829 2663 2835 2677
rect 3012 2677 3068 2683
rect 3108 2677 3132 2683
rect 3149 2677 3180 2683
rect 2740 2657 2835 2663
rect 3149 2663 3155 2677
rect 3677 2683 3683 2697
rect 3732 2697 3788 2703
rect 3812 2697 4019 2703
rect 4013 2684 4019 2697
rect 4052 2697 4108 2703
rect 4276 2697 4348 2703
rect 4356 2697 4476 2703
rect 4500 2697 4780 2703
rect 4852 2697 5020 2703
rect 5252 2697 5708 2703
rect 5716 2697 5756 2703
rect 5885 2703 5891 2717
rect 5956 2717 6076 2723
rect 6132 2717 6227 2723
rect 5812 2697 5891 2703
rect 5908 2697 6108 2703
rect 6164 2697 6204 2703
rect 3677 2677 3772 2683
rect 3812 2677 3836 2683
rect 3853 2677 3916 2683
rect 2852 2657 3155 2663
rect 3284 2657 3308 2663
rect 3364 2657 3468 2663
rect 3668 2657 3676 2663
rect 3700 2657 3724 2663
rect 3853 2663 3859 2677
rect 3933 2677 4003 2683
rect 3764 2657 3859 2663
rect 3876 2657 3884 2663
rect 3933 2663 3939 2677
rect 3924 2657 3939 2663
rect 3956 2657 3980 2663
rect 3997 2663 4003 2677
rect 4036 2677 4163 2683
rect 3997 2657 4012 2663
rect 4020 2657 4108 2663
rect 4157 2663 4163 2677
rect 4180 2677 4492 2683
rect 4516 2677 4588 2683
rect 4868 2677 4892 2683
rect 4900 2677 4908 2683
rect 5236 2677 5772 2683
rect 5780 2677 5868 2683
rect 5876 2677 6188 2683
rect 6221 2664 6227 2717
rect 4157 2657 4316 2663
rect 4324 2657 4396 2663
rect 4452 2657 4652 2663
rect 4660 2657 4764 2663
rect 4772 2657 4876 2663
rect 4884 2657 4972 2663
rect 5076 2657 5196 2663
rect 5204 2657 5308 2663
rect 5492 2657 5740 2663
rect 5812 2657 5932 2663
rect 5988 2657 6012 2663
rect 6036 2657 6092 2663
rect 6132 2657 6188 2663
rect 2269 2637 2364 2643
rect 2420 2637 2508 2643
rect 2532 2637 2700 2643
rect 2756 2637 2908 2643
rect 2916 2637 3100 2643
rect 3124 2637 3276 2643
rect 3284 2637 3292 2643
rect 3316 2637 3532 2643
rect 3620 2637 5548 2643
rect 5556 2637 5612 2643
rect 5620 2637 5932 2643
rect 5972 2637 6044 2643
rect 6084 2637 6124 2643
rect 6132 2637 6156 2643
rect 260 2617 284 2623
rect 452 2617 460 2623
rect 516 2617 620 2623
rect 932 2617 1068 2623
rect 1076 2617 1132 2623
rect 1172 2617 1820 2623
rect 1844 2617 1868 2623
rect 1956 2617 2028 2623
rect 2148 2617 2220 2623
rect 2260 2617 2300 2623
rect 2388 2617 2636 2623
rect 2660 2617 2732 2623
rect 2772 2617 2876 2623
rect 2893 2617 2988 2623
rect 308 2597 348 2603
rect 356 2597 716 2603
rect 852 2597 988 2603
rect 1012 2597 2220 2603
rect 2356 2597 2620 2603
rect 2708 2597 2796 2603
rect 2893 2603 2899 2617
rect 3060 2617 3084 2623
rect 3188 2617 3452 2623
rect 3476 2617 3500 2623
rect 3524 2617 3747 2623
rect 3112 2614 3160 2616
rect 3112 2606 3113 2614
rect 3122 2606 3123 2614
rect 3158 2606 3160 2614
rect 3112 2604 3160 2606
rect 2804 2597 2899 2603
rect 2964 2597 2988 2603
rect 3044 2597 3068 2603
rect 3204 2597 3404 2603
rect 3444 2597 3468 2603
rect 3492 2597 3500 2603
rect 3572 2597 3628 2603
rect 3668 2597 3724 2603
rect 3741 2603 3747 2617
rect 3764 2617 3916 2623
rect 4004 2617 4172 2623
rect 4244 2617 4508 2623
rect 5300 2617 5324 2623
rect 5348 2617 5500 2623
rect 5508 2617 5580 2623
rect 5748 2617 5788 2623
rect 5812 2617 5852 2623
rect 5908 2617 5996 2623
rect 3741 2597 3804 2603
rect 3828 2597 3852 2603
rect 3860 2597 4236 2603
rect 4253 2597 4396 2603
rect 100 2577 108 2583
rect 324 2577 332 2583
rect 340 2577 508 2583
rect 612 2577 1100 2583
rect 1124 2577 1180 2583
rect 1396 2577 1484 2583
rect 1572 2577 1964 2583
rect 2020 2577 2044 2583
rect 2068 2577 2412 2583
rect 2484 2577 2796 2583
rect 2884 2577 3196 2583
rect 3236 2577 3260 2583
rect 3316 2577 3484 2583
rect 3508 2577 3564 2583
rect 3604 2577 3996 2583
rect 4052 2577 4172 2583
rect 4253 2583 4259 2597
rect 4436 2597 4476 2603
rect 4596 2597 4764 2603
rect 5396 2597 5708 2603
rect 5716 2597 5932 2603
rect 6020 2597 6124 2603
rect 6132 2597 6156 2603
rect 6237 2597 6300 2603
rect 4212 2577 4259 2583
rect 4372 2577 4620 2583
rect 4660 2577 4716 2583
rect 4948 2577 4988 2583
rect 4996 2577 5020 2583
rect 5492 2577 6003 2583
rect 5997 2564 6003 2577
rect 6036 2577 6124 2583
rect 6237 2583 6243 2597
rect 6141 2577 6243 2583
rect 52 2557 204 2563
rect 500 2557 556 2563
rect 628 2557 716 2563
rect 756 2557 940 2563
rect 948 2557 972 2563
rect 1220 2557 1308 2563
rect 1556 2557 1564 2563
rect 1604 2557 1660 2563
rect 1700 2557 1852 2563
rect 1876 2557 1900 2563
rect 1924 2557 1996 2563
rect 2020 2557 2092 2563
rect 2100 2557 2172 2563
rect 2196 2557 2300 2563
rect 2452 2557 2524 2563
rect 2541 2557 2588 2563
rect 20 2537 44 2543
rect 100 2537 140 2543
rect 308 2537 364 2543
rect 468 2537 524 2543
rect 580 2537 620 2543
rect 660 2537 844 2543
rect 884 2537 972 2543
rect 996 2537 1292 2543
rect 1332 2537 1356 2543
rect 1412 2537 1676 2543
rect 1684 2537 1756 2543
rect 1828 2537 1884 2543
rect 1988 2537 2012 2543
rect 2036 2537 2060 2543
rect 2196 2537 2316 2543
rect 2340 2537 2396 2543
rect 2420 2537 2476 2543
rect 2541 2543 2547 2557
rect 2644 2557 2716 2563
rect 2740 2557 2844 2563
rect 2964 2557 3052 2563
rect 3076 2557 3180 2563
rect 3204 2557 3244 2563
rect 3332 2557 3372 2563
rect 3412 2557 3436 2563
rect 3460 2557 3692 2563
rect 3812 2557 3820 2563
rect 3844 2557 3980 2563
rect 4004 2557 4060 2563
rect 4116 2557 4284 2563
rect 4484 2557 4508 2563
rect 4516 2557 4652 2563
rect 5588 2557 5772 2563
rect 6141 2563 6147 2577
rect 6084 2557 6147 2563
rect 6164 2557 6188 2563
rect 2500 2537 2547 2543
rect 2564 2537 2604 2543
rect 2708 2537 2764 2543
rect 2836 2537 2892 2543
rect 2948 2537 3052 2543
rect 3092 2537 3244 2543
rect 3300 2537 3324 2543
rect 3380 2537 3500 2543
rect 3540 2537 3580 2543
rect 3796 2537 3916 2543
rect 3940 2537 4140 2543
rect 4148 2537 4524 2543
rect 4740 2537 4860 2543
rect 4932 2537 5132 2543
rect 5268 2537 5324 2543
rect 5364 2537 5436 2543
rect 5460 2537 5644 2543
rect 5764 2537 5836 2543
rect 5972 2537 6035 2543
rect 20 2517 28 2523
rect 132 2517 284 2523
rect 308 2517 396 2523
rect 436 2517 540 2523
rect 580 2517 732 2523
rect 820 2517 1164 2523
rect 1204 2517 1260 2523
rect 1284 2517 1356 2523
rect 1396 2517 1772 2523
rect 1780 2517 2092 2523
rect 2132 2517 2524 2523
rect 2644 2517 3820 2523
rect 3876 2517 3916 2523
rect 3972 2517 4012 2523
rect 4084 2517 4092 2523
rect 4116 2517 4140 2523
rect 4180 2517 4300 2523
rect 4372 2517 4460 2523
rect 4525 2523 4531 2536
rect 6029 2524 6035 2537
rect 6116 2537 6156 2543
rect 6173 2537 6252 2543
rect 4525 2517 5692 2523
rect 5700 2517 5804 2523
rect 5844 2517 5964 2523
rect 6173 2523 6179 2537
rect 6068 2517 6179 2523
rect 548 2497 556 2503
rect 596 2497 652 2503
rect 724 2497 780 2503
rect 884 2497 1020 2503
rect 1108 2497 1148 2503
rect 1204 2497 1244 2503
rect 1332 2497 1948 2503
rect 2004 2497 2060 2503
rect 2077 2497 2156 2503
rect 500 2477 540 2483
rect 548 2477 684 2483
rect 756 2477 988 2483
rect 1076 2477 1148 2483
rect 1172 2477 1388 2483
rect 1412 2477 1443 2483
rect 660 2457 684 2463
rect 724 2457 876 2463
rect 900 2457 1132 2463
rect 1316 2457 1340 2463
rect 1380 2457 1420 2463
rect 772 2437 1420 2443
rect 1437 2443 1443 2477
rect 1460 2477 1500 2483
rect 1508 2477 1516 2483
rect 1540 2477 1628 2483
rect 1684 2477 1708 2483
rect 1860 2477 2012 2483
rect 2077 2483 2083 2497
rect 2308 2497 2332 2503
rect 2436 2497 2620 2503
rect 2852 2497 2892 2503
rect 2996 2497 3084 2503
rect 3108 2497 3404 2503
rect 3444 2497 3683 2503
rect 2397 2484 2403 2496
rect 2036 2477 2083 2483
rect 2100 2477 2380 2483
rect 2420 2477 2716 2483
rect 2740 2477 2780 2483
rect 2788 2477 2860 2483
rect 2868 2477 2908 2483
rect 2932 2477 3084 2483
rect 3140 2477 3212 2483
rect 3236 2477 3468 2483
rect 3492 2477 3564 2483
rect 3677 2483 3683 2497
rect 3700 2497 3836 2503
rect 3924 2497 3948 2503
rect 3988 2497 4044 2503
rect 4116 2497 4140 2503
rect 4180 2497 4252 2503
rect 4276 2497 4332 2503
rect 4436 2497 4540 2503
rect 4900 2497 4956 2503
rect 5108 2497 5212 2503
rect 5300 2497 5516 2503
rect 5524 2497 5628 2503
rect 5716 2497 5788 2503
rect 5812 2497 5916 2503
rect 6052 2497 6156 2503
rect 3677 2477 3756 2483
rect 3796 2477 3884 2483
rect 3892 2477 4476 2483
rect 5428 2477 5436 2483
rect 5764 2477 5772 2483
rect 6205 2483 6211 2516
rect 6269 2484 6275 2576
rect 6052 2477 6211 2483
rect 1460 2457 3100 2463
rect 3220 2457 3276 2463
rect 3293 2457 3372 2463
rect 1437 2437 1452 2443
rect 1524 2437 1724 2443
rect 1764 2437 1852 2443
rect 1892 2437 2092 2443
rect 2372 2437 2812 2443
rect 2836 2437 2876 2443
rect 2932 2437 2972 2443
rect 2996 2437 3020 2443
rect 3293 2443 3299 2457
rect 3380 2457 3427 2463
rect 3421 2444 3427 2457
rect 3444 2457 3692 2463
rect 3709 2457 3868 2463
rect 3044 2437 3299 2443
rect 3316 2437 3388 2443
rect 3460 2437 3532 2443
rect 3588 2437 3628 2443
rect 3709 2443 3715 2457
rect 3892 2457 4364 2463
rect 5940 2457 6108 2463
rect 3684 2437 3715 2443
rect 3860 2437 3932 2443
rect 3956 2437 3980 2443
rect 4036 2437 4092 2443
rect 4148 2437 4236 2443
rect 4276 2437 4332 2443
rect 4340 2437 4444 2443
rect 4452 2437 4572 2443
rect 4580 2437 4620 2443
rect 4628 2437 4748 2443
rect 5556 2437 5612 2443
rect 5620 2437 5692 2443
rect 5700 2437 5724 2443
rect 5732 2437 5740 2443
rect 6036 2437 6092 2443
rect 6100 2437 6220 2443
rect 676 2417 684 2423
rect 772 2417 828 2423
rect 836 2417 908 2423
rect 948 2417 1452 2423
rect 1668 2417 1708 2423
rect 1940 2417 2060 2423
rect 2084 2417 2956 2423
rect 3028 2417 3228 2423
rect 3252 2417 3660 2423
rect 3748 2417 3756 2423
rect 3764 2417 4284 2423
rect 4308 2417 4524 2423
rect 5732 2417 5900 2423
rect 1576 2414 1624 2416
rect 1576 2406 1577 2414
rect 1586 2406 1587 2414
rect 1622 2406 1624 2414
rect 1576 2404 1624 2406
rect 4664 2414 4712 2416
rect 4664 2406 4665 2414
rect 4674 2406 4675 2414
rect 4710 2406 4712 2414
rect 4664 2404 4712 2406
rect 468 2397 476 2403
rect 644 2397 796 2403
rect 804 2397 1404 2403
rect 1428 2397 1484 2403
rect 1652 2397 1836 2403
rect 2100 2397 2108 2403
rect 2260 2397 2268 2403
rect 2324 2397 2636 2403
rect 2724 2397 3180 2403
rect 3213 2397 3324 2403
rect 84 2377 140 2383
rect 148 2377 764 2383
rect 820 2377 844 2383
rect 852 2377 1516 2383
rect 1540 2377 1820 2383
rect 1837 2377 1884 2383
rect 420 2357 508 2363
rect 516 2357 620 2363
rect 628 2357 668 2363
rect 676 2357 748 2363
rect 788 2357 828 2363
rect 836 2357 924 2363
rect 932 2357 1500 2363
rect 1524 2357 1580 2363
rect 1652 2357 1724 2363
rect 1837 2363 1843 2377
rect 1956 2377 2380 2383
rect 2404 2377 2476 2383
rect 2516 2377 2604 2383
rect 2628 2377 2668 2383
rect 2740 2377 2828 2383
rect 2852 2377 2860 2383
rect 2868 2377 2924 2383
rect 2932 2377 2988 2383
rect 3213 2383 3219 2397
rect 3332 2397 3468 2403
rect 3476 2397 3916 2403
rect 4004 2397 4028 2403
rect 4052 2397 4396 2403
rect 4436 2397 4476 2403
rect 5076 2397 5228 2403
rect 5812 2397 6275 2403
rect 3060 2377 3219 2383
rect 3236 2377 3292 2383
rect 3316 2377 3564 2383
rect 3620 2377 3836 2383
rect 3908 2377 4124 2383
rect 4132 2377 4252 2383
rect 4276 2377 4284 2383
rect 4324 2377 4668 2383
rect 4772 2377 5772 2383
rect 6148 2377 6188 2383
rect 1796 2357 1843 2363
rect 1860 2357 1868 2363
rect 1876 2357 2028 2363
rect 2068 2357 2124 2363
rect 2228 2357 2364 2363
rect 2420 2357 2636 2363
rect 2660 2357 2796 2363
rect 2804 2357 3052 2363
rect 3060 2357 3644 2363
rect 3652 2357 5068 2363
rect 5988 2357 6060 2363
rect 356 2337 428 2343
rect 532 2337 652 2343
rect 692 2337 940 2343
rect 1012 2337 1196 2343
rect 1300 2337 1388 2343
rect 1460 2337 1907 2343
rect 1901 2324 1907 2337
rect 1972 2337 2124 2343
rect 2372 2337 2428 2343
rect 2468 2337 2556 2343
rect 2596 2337 2684 2343
rect 2884 2337 2892 2343
rect 2900 2337 2940 2343
rect 2948 2337 3084 2343
rect 3101 2337 3340 2343
rect 2221 2324 2227 2336
rect 308 2317 332 2323
rect 340 2317 428 2323
rect 436 2317 524 2323
rect 548 2317 732 2323
rect 788 2317 844 2323
rect 868 2317 892 2323
rect 1044 2317 1324 2323
rect 1332 2317 1388 2323
rect 1412 2317 1484 2323
rect 1524 2317 1644 2323
rect 1716 2317 1788 2323
rect 1796 2317 1884 2323
rect 1940 2317 2220 2323
rect 2244 2317 2300 2323
rect 2436 2317 2492 2323
rect 2580 2317 2764 2323
rect 3101 2323 3107 2337
rect 3396 2337 3884 2343
rect 3924 2337 4156 2343
rect 4196 2337 4332 2343
rect 4356 2337 4380 2343
rect 4420 2337 4476 2343
rect 4532 2337 4588 2343
rect 5252 2337 5324 2343
rect 5684 2337 5772 2343
rect 6052 2337 6060 2343
rect 6212 2337 6252 2343
rect 6269 2343 6275 2397
rect 6269 2337 6291 2343
rect 6285 2324 6291 2337
rect 2996 2317 3107 2323
rect 3124 2317 3868 2323
rect 3876 2317 4124 2323
rect 4132 2317 4748 2323
rect 4756 2317 4988 2323
rect 5620 2317 5644 2323
rect 6164 2317 6259 2323
rect -19 2297 12 2303
rect 196 2297 524 2303
rect 644 2297 892 2303
rect 916 2297 956 2303
rect 980 2297 1116 2303
rect 1220 2297 2076 2303
rect 2100 2297 2156 2303
rect 2260 2297 2371 2303
rect 68 2277 300 2283
rect 388 2277 540 2283
rect 573 2283 579 2296
rect 564 2277 643 2283
rect 148 2257 332 2263
rect 580 2257 620 2263
rect 637 2263 643 2277
rect 660 2277 684 2283
rect 788 2277 940 2283
rect 980 2277 1068 2283
rect 1172 2277 1276 2283
rect 1332 2277 1356 2283
rect 1428 2277 1548 2283
rect 1700 2277 1740 2283
rect 1764 2277 1820 2283
rect 1828 2277 1964 2283
rect 1988 2277 2115 2283
rect 637 2257 1020 2263
rect 1444 2257 1660 2263
rect 1684 2257 1724 2263
rect 1796 2257 1964 2263
rect 1972 2257 2092 2263
rect 2109 2263 2115 2277
rect 2180 2277 2236 2283
rect 2253 2277 2316 2283
rect 2109 2257 2172 2263
rect 2253 2263 2259 2277
rect 2365 2283 2371 2297
rect 2388 2297 2476 2303
rect 2548 2297 2588 2303
rect 2612 2297 2675 2303
rect 2365 2277 2492 2283
rect 2500 2277 2540 2283
rect 2564 2277 2572 2283
rect 2596 2280 2604 2283
rect 2596 2277 2611 2280
rect 2644 2277 2652 2283
rect 2669 2283 2675 2297
rect 2756 2297 2764 2303
rect 2781 2303 2787 2316
rect 2781 2297 3004 2303
rect 3028 2297 3100 2303
rect 3124 2297 3532 2303
rect 3620 2297 3628 2303
rect 3796 2297 3932 2303
rect 4068 2297 4204 2303
rect 4212 2297 4316 2303
rect 4324 2297 4492 2303
rect 4500 2297 5068 2303
rect 5076 2297 5100 2303
rect 5284 2297 5372 2303
rect 5588 2297 5644 2303
rect 5748 2297 5804 2303
rect 5677 2284 5683 2296
rect 2669 2277 2844 2283
rect 2868 2277 2876 2283
rect 2916 2277 3036 2283
rect 3060 2277 3244 2283
rect 3268 2277 3372 2283
rect 3485 2277 3516 2283
rect 2196 2257 2259 2263
rect 2276 2257 2316 2263
rect 2340 2257 2444 2263
rect 2516 2257 2524 2263
rect 2532 2257 2588 2263
rect 2605 2260 2668 2263
rect 429 2244 435 2256
rect 2612 2257 2668 2260
rect 2692 2257 2748 2263
rect 2772 2257 2828 2263
rect 2916 2257 2924 2263
rect 2964 2257 3020 2263
rect 3069 2257 3116 2263
rect 532 2237 780 2243
rect 804 2237 1452 2243
rect 1460 2237 1836 2243
rect 1844 2237 1852 2243
rect 3069 2243 3075 2257
rect 3188 2257 3228 2263
rect 3284 2257 3436 2263
rect 3485 2263 3491 2277
rect 3540 2277 3596 2283
rect 3636 2277 3692 2283
rect 3764 2277 3875 2283
rect 3693 2264 3699 2276
rect 3476 2257 3491 2263
rect 3501 2257 3548 2263
rect 1876 2237 3075 2243
rect 3108 2237 3212 2243
rect 3229 2237 3308 2243
rect 692 2217 796 2223
rect 820 2217 844 2223
rect 1044 2217 1804 2223
rect 1924 2217 2156 2223
rect 2164 2217 2732 2223
rect 2804 2217 2924 2223
rect 2948 2217 2972 2223
rect 3012 2217 3084 2223
rect 3229 2223 3235 2237
rect 3348 2237 3420 2243
rect 3428 2237 3452 2243
rect 3501 2243 3507 2257
rect 3604 2257 3644 2263
rect 3732 2257 3788 2263
rect 3828 2257 3852 2263
rect 3869 2263 3875 2277
rect 3892 2277 3996 2283
rect 4148 2277 4156 2283
rect 4244 2277 4348 2283
rect 4388 2277 4460 2283
rect 4516 2277 4636 2283
rect 4644 2277 4652 2283
rect 4724 2277 4892 2283
rect 5428 2277 5516 2283
rect 5844 2277 5916 2283
rect 5940 2277 5948 2283
rect 6004 2277 6156 2283
rect 3869 2257 3900 2263
rect 3924 2257 4140 2263
rect 4148 2257 4236 2263
rect 4292 2257 4364 2263
rect 4436 2257 4812 2263
rect 4820 2257 4860 2263
rect 5700 2257 5804 2263
rect 6052 2257 6236 2263
rect 3492 2237 3507 2243
rect 3524 2237 3628 2243
rect 3668 2237 3724 2243
rect 3748 2237 4108 2243
rect 4292 2237 4444 2243
rect 4468 2237 4476 2243
rect 4484 2237 4556 2243
rect 4580 2237 4636 2243
rect 4660 2237 4796 2243
rect 4804 2237 4828 2243
rect 4868 2237 5004 2243
rect 5044 2237 5804 2243
rect 5956 2237 6012 2243
rect 6253 2243 6259 2317
rect 6228 2237 6259 2243
rect 3220 2217 3235 2223
rect 3316 2217 3372 2223
rect 3476 2217 3692 2223
rect 3764 2217 5164 2223
rect 5684 2217 6252 2223
rect 3112 2214 3160 2216
rect 3112 2206 3113 2214
rect 3122 2206 3123 2214
rect 3158 2206 3160 2214
rect 3112 2204 3160 2206
rect 372 2197 428 2203
rect 660 2197 748 2203
rect 820 2197 1068 2203
rect 1092 2197 1212 2203
rect 1268 2197 1868 2203
rect 1892 2197 2028 2203
rect 2036 2197 2060 2203
rect 2116 2197 2188 2203
rect 2276 2197 2348 2203
rect 2365 2197 2396 2203
rect 500 2177 1260 2183
rect 1332 2177 1404 2183
rect 1428 2177 1740 2183
rect 1812 2177 1836 2183
rect 1940 2177 1948 2183
rect 1956 2177 2044 2183
rect 2077 2177 2252 2183
rect 148 2157 204 2163
rect 260 2157 300 2163
rect 356 2157 428 2163
rect 436 2157 652 2163
rect 820 2157 844 2163
rect 1012 2157 1020 2163
rect 132 2137 524 2143
rect 596 2137 924 2143
rect 941 2137 1020 2143
rect 180 2117 316 2123
rect 468 2117 620 2123
rect 941 2123 947 2137
rect 1044 2137 1116 2143
rect 1156 2137 1180 2143
rect 1268 2137 1372 2143
rect 1405 2143 1411 2176
rect 1460 2157 1500 2163
rect 1716 2157 1724 2163
rect 1780 2157 1868 2163
rect 2077 2163 2083 2177
rect 2365 2183 2371 2197
rect 2420 2197 2460 2203
rect 2484 2197 2668 2203
rect 2772 2197 3052 2203
rect 3188 2197 3468 2203
rect 3476 2197 3884 2203
rect 3988 2197 4300 2203
rect 4372 2197 4476 2203
rect 4564 2197 4588 2203
rect 4612 2197 4780 2203
rect 5028 2197 5036 2203
rect 5684 2197 5708 2203
rect 5716 2197 5820 2203
rect 5876 2197 6028 2203
rect 6084 2197 6115 2203
rect 2292 2177 2371 2183
rect 2452 2177 2492 2183
rect 2564 2177 2684 2183
rect 2692 2177 2716 2183
rect 2772 2177 2860 2183
rect 2884 2177 3091 2183
rect 1972 2157 2083 2163
rect 2100 2157 2124 2163
rect 2141 2157 2332 2163
rect 1405 2137 1564 2143
rect 1661 2137 1676 2143
rect 660 2117 947 2123
rect 980 2117 1084 2123
rect 1140 2117 1164 2123
rect 1204 2117 1228 2123
rect 1236 2117 1324 2123
rect 1661 2123 1667 2137
rect 1684 2137 1708 2143
rect 1732 2137 1932 2143
rect 2004 2137 2012 2143
rect 2141 2143 2147 2157
rect 2356 2157 2460 2163
rect 2468 2157 2476 2163
rect 2500 2157 2540 2163
rect 2612 2157 2636 2163
rect 2676 2157 2796 2163
rect 2820 2157 2844 2163
rect 2884 2157 3068 2163
rect 3085 2163 3091 2177
rect 3108 2177 3388 2183
rect 3412 2177 3516 2183
rect 3572 2177 3612 2183
rect 3629 2177 3900 2183
rect 3085 2157 3308 2163
rect 3380 2157 3484 2163
rect 3629 2163 3635 2177
rect 3924 2177 4172 2183
rect 4244 2177 4252 2183
rect 4260 2177 4380 2183
rect 4436 2177 4620 2183
rect 4644 2177 4812 2183
rect 4884 2177 5132 2183
rect 5188 2177 5804 2183
rect 5812 2177 5836 2183
rect 5844 2177 6092 2183
rect 3540 2157 3635 2163
rect 3652 2157 3820 2163
rect 3844 2157 3907 2163
rect 2020 2137 2147 2143
rect 2164 2137 2572 2143
rect 2756 2137 2988 2143
rect 3092 2137 3228 2143
rect 3236 2137 3395 2143
rect 1332 2117 1667 2123
rect 1684 2117 1708 2123
rect 1812 2117 1884 2123
rect 1933 2117 2956 2123
rect 84 2097 204 2103
rect 308 2097 364 2103
rect 372 2097 556 2103
rect 580 2097 716 2103
rect 740 2097 892 2103
rect 1005 2097 1228 2103
rect 484 2077 556 2083
rect 1005 2083 1011 2097
rect 1604 2097 1660 2103
rect 1933 2103 1939 2117
rect 3389 2123 3395 2137
rect 3428 2137 3516 2143
rect 3540 2137 3756 2143
rect 3860 2137 3868 2143
rect 3901 2143 3907 2157
rect 3924 2157 4099 2163
rect 3901 2137 3932 2143
rect 4093 2143 4099 2157
rect 4132 2157 4204 2163
rect 4276 2157 4492 2163
rect 4596 2157 5084 2163
rect 5828 2157 5852 2163
rect 6109 2163 6115 2197
rect 6148 2197 6188 2203
rect 6100 2157 6115 2163
rect 4269 2144 4275 2156
rect 4093 2137 4204 2143
rect 4340 2137 4396 2143
rect 4429 2137 4460 2143
rect 2980 2117 3379 2123
rect 3389 2117 3491 2123
rect 1796 2097 1939 2103
rect 2004 2097 2012 2103
rect 2068 2097 2108 2103
rect 2180 2097 2204 2103
rect 2228 2097 2236 2103
rect 2340 2097 2476 2103
rect 2516 2097 2540 2103
rect 2580 2097 2716 2103
rect 2740 2097 2780 2103
rect 2804 2097 2988 2103
rect 3012 2097 3132 2103
rect 3140 2097 3148 2103
rect 3156 2097 3244 2103
rect 3332 2097 3356 2103
rect 3373 2103 3379 2117
rect 3373 2097 3404 2103
rect 3485 2103 3491 2117
rect 3508 2117 3564 2123
rect 3597 2117 3628 2123
rect 3597 2103 3603 2117
rect 3700 2117 3724 2123
rect 3796 2117 3852 2123
rect 3876 2117 4364 2123
rect 4429 2123 4435 2137
rect 4484 2137 4716 2143
rect 4724 2137 5004 2143
rect 5060 2137 5116 2143
rect 5124 2137 5212 2143
rect 5364 2137 5500 2143
rect 5508 2137 5676 2143
rect 6036 2137 6076 2143
rect 4372 2117 4435 2123
rect 4452 2117 4556 2123
rect 4564 2117 4588 2123
rect 4708 2117 4732 2123
rect 4836 2117 4844 2123
rect 4868 2117 4940 2123
rect 5156 2117 5260 2123
rect 5332 2117 5356 2123
rect 5428 2117 5468 2123
rect 5828 2117 5852 2123
rect 5876 2117 6012 2123
rect 5037 2104 5043 2116
rect 3485 2097 3603 2103
rect 3620 2097 3676 2103
rect 3780 2097 3852 2103
rect 3940 2097 3964 2103
rect 3988 2097 4060 2103
rect 4084 2097 4108 2103
rect 4260 2097 4284 2103
rect 4308 2097 4380 2103
rect 4404 2097 5004 2103
rect 5140 2097 5916 2103
rect 596 2077 1011 2083
rect 1028 2077 1068 2083
rect 1156 2077 1164 2083
rect 1172 2077 1196 2083
rect 1220 2077 1372 2083
rect 1396 2077 1532 2083
rect 1757 2083 1763 2096
rect 6269 2084 6275 2176
rect 1757 2077 1804 2083
rect 1812 2077 1900 2083
rect 1924 2077 1980 2083
rect 2004 2077 2172 2083
rect 2180 2077 2780 2083
rect 2788 2077 2860 2083
rect 2868 2077 2940 2083
rect 2996 2077 3020 2083
rect 3028 2077 3164 2083
rect 3188 2077 3244 2083
rect 3252 2077 3500 2083
rect 3508 2077 3660 2083
rect 3668 2077 4316 2083
rect 4340 2077 4588 2083
rect 4596 2077 4620 2083
rect 4756 2077 5324 2083
rect 5844 2077 6028 2083
rect 6036 2077 6108 2083
rect 6116 2077 6156 2083
rect 436 2057 492 2063
rect 564 2057 604 2063
rect 772 2057 988 2063
rect 996 2057 1324 2063
rect 1652 2057 1692 2063
rect 1780 2057 2812 2063
rect 2820 2057 2860 2063
rect 2884 2057 2956 2063
rect 2996 2057 3020 2063
rect 3044 2057 3340 2063
rect 3364 2057 3916 2063
rect 3956 2057 3996 2063
rect 4020 2057 4108 2063
rect 4164 2057 4236 2063
rect 4420 2057 4460 2063
rect 4516 2057 4604 2063
rect 4644 2057 4876 2063
rect 5044 2057 5100 2063
rect 5332 2057 5388 2063
rect 6068 2057 6092 2063
rect 884 2037 2364 2043
rect 2548 2037 2604 2043
rect 2644 2037 4028 2043
rect 4052 2037 4172 2043
rect 4244 2037 4268 2043
rect 4372 2037 4764 2043
rect 4788 2037 4796 2043
rect 4852 2037 5196 2043
rect 5613 2024 5619 2036
rect 404 2017 476 2023
rect 516 2017 780 2023
rect 852 2017 892 2023
rect 900 2017 908 2023
rect 1076 2017 1212 2023
rect 1348 2017 1388 2023
rect 1412 2017 1468 2023
rect 1668 2017 1836 2023
rect 1844 2017 2332 2023
rect 2356 2017 2380 2023
rect 2404 2017 2476 2023
rect 2500 2017 2540 2023
rect 2612 2017 2620 2023
rect 2644 2017 2652 2023
rect 2724 2017 2764 2023
rect 2820 2017 2876 2023
rect 2900 2017 2972 2023
rect 2980 2017 3180 2023
rect 3204 2017 3235 2023
rect 1576 2014 1624 2016
rect 1576 2006 1577 2014
rect 1586 2006 1587 2014
rect 1622 2006 1624 2014
rect 1576 2004 1624 2006
rect 20 1997 412 2003
rect 420 1997 476 2003
rect 484 1997 972 2003
rect 980 1997 1068 2003
rect 1092 1997 1132 2003
rect 1156 1997 1196 2003
rect 1252 1997 1276 2003
rect 1284 1997 1340 2003
rect 1380 1997 1404 2003
rect 1492 1997 1516 2003
rect 1668 1997 1676 2003
rect 1716 1997 1756 2003
rect 1812 1997 1964 2003
rect 1972 1997 2220 2003
rect 2228 1997 2508 2003
rect 2628 1997 2716 2003
rect 2900 1997 3212 2003
rect 3229 2003 3235 2017
rect 3268 2017 3292 2023
rect 3300 2017 3628 2023
rect 3668 2017 4636 2023
rect 4820 2017 5020 2023
rect 5780 2017 6028 2023
rect 6052 2017 6092 2023
rect 6164 2017 6188 2023
rect 4664 2014 4712 2016
rect 4664 2006 4665 2014
rect 4674 2006 4675 2014
rect 4710 2006 4712 2014
rect 4664 2004 4712 2006
rect 3229 1997 3276 2003
rect 3325 1997 3340 2003
rect 356 1977 492 1983
rect 548 1977 620 1983
rect 644 1977 668 1983
rect 916 1977 1036 1983
rect 1044 1977 1804 1983
rect 1844 1977 1868 1983
rect 1956 1977 1980 1983
rect 2004 1977 2044 1983
rect 2100 1977 2140 1983
rect 2148 1977 2172 1983
rect 2196 1977 2252 1983
rect 2356 1977 2387 1983
rect 404 1957 428 1963
rect 500 1957 972 1963
rect 989 1957 1068 1963
rect 452 1937 556 1943
rect 564 1937 572 1943
rect 660 1937 732 1943
rect 989 1943 995 1957
rect 1092 1957 1244 1963
rect 1252 1957 1276 1963
rect 1284 1957 1324 1963
rect 1332 1957 1388 1963
rect 1428 1957 1667 1963
rect 788 1937 995 1943
rect 1028 1937 1164 1943
rect 1172 1937 1484 1943
rect 1492 1937 1644 1943
rect 1661 1943 1667 1957
rect 1684 1957 1868 1963
rect 1892 1957 2124 1963
rect 2228 1957 2252 1963
rect 2381 1963 2387 1977
rect 2452 1977 2476 1983
rect 2548 1977 2812 1983
rect 2852 1977 3100 1983
rect 3188 1977 3212 1983
rect 3325 1983 3331 1997
rect 3412 1997 3532 2003
rect 3556 1997 3580 2003
rect 3604 1997 3660 2003
rect 3684 1997 3779 2003
rect 3220 1977 3331 1983
rect 3348 1977 3756 1983
rect 3773 1983 3779 1997
rect 3812 1997 3980 2003
rect 4052 1997 4140 2003
rect 4164 1997 4611 2003
rect 3773 1977 3820 1983
rect 3956 1977 3964 1983
rect 4004 1977 4428 1983
rect 4605 1983 4611 1997
rect 5012 1997 6092 2003
rect 6196 1997 6300 2003
rect 4605 1977 4652 1983
rect 4708 1977 4732 1983
rect 4996 1977 5420 1983
rect 5716 1977 5804 1983
rect 6164 1977 6195 1983
rect 6189 1964 6195 1977
rect 2381 1957 2588 1963
rect 2596 1957 2748 1963
rect 2868 1957 2892 1963
rect 2932 1957 3020 1963
rect 3108 1957 3276 1963
rect 3316 1957 3612 1963
rect 3620 1957 4044 1963
rect 4068 1957 4092 1963
rect 4308 1957 4348 1963
rect 4404 1957 4508 1963
rect 4596 1957 5164 1963
rect 5748 1957 5932 1963
rect 5988 1957 6012 1963
rect 6100 1957 6156 1963
rect 6212 1957 6268 1963
rect 1661 1937 1900 1943
rect 1940 1937 2012 1943
rect 2077 1937 2124 1943
rect 148 1917 284 1923
rect 436 1917 588 1923
rect 596 1917 620 1923
rect 628 1917 828 1923
rect 836 1917 1132 1923
rect 1188 1917 1244 1923
rect 1300 1917 1324 1923
rect 1501 1917 1603 1923
rect 116 1897 204 1903
rect 244 1897 284 1903
rect 372 1897 380 1903
rect 388 1897 748 1903
rect 900 1897 1100 1903
rect 1501 1903 1507 1917
rect 1149 1897 1507 1903
rect 1597 1903 1603 1917
rect 1620 1917 1708 1923
rect 1732 1917 1740 1923
rect 2077 1923 2083 1937
rect 2164 1937 2220 1943
rect 2340 1937 2540 1943
rect 2948 1937 3212 1943
rect 3268 1937 3356 1943
rect 3428 1937 3660 1943
rect 3684 1937 3708 1943
rect 3748 1937 3852 1943
rect 3860 1937 4604 1943
rect 4644 1937 4732 1943
rect 4740 1937 4844 1943
rect 4852 1937 4876 1943
rect 5060 1937 5084 1943
rect 5204 1937 5228 1943
rect 5252 1937 5340 1943
rect 5364 1937 5404 1943
rect 5572 1937 5596 1943
rect 5748 1937 6108 1943
rect 6132 1937 6156 1943
rect 1764 1917 2083 1923
rect 2164 1917 2172 1923
rect 2244 1917 2412 1923
rect 2548 1917 2620 1923
rect 2644 1920 2924 1923
rect 2644 1917 2931 1920
rect 2964 1917 3100 1923
rect 3124 1917 3244 1923
rect 3316 1917 3340 1923
rect 3364 1917 3388 1923
rect 3396 1917 3459 1923
rect 1597 1897 1676 1903
rect 1149 1884 1155 1897
rect 1732 1897 1804 1903
rect 1876 1897 1900 1903
rect 1940 1897 1964 1903
rect 1988 1897 2028 1903
rect 2068 1897 2140 1903
rect 2196 1897 2828 1903
rect 2932 1897 3036 1903
rect 3092 1897 3356 1903
rect 3396 1897 3436 1903
rect 3453 1903 3459 1917
rect 3476 1917 3516 1923
rect 3540 1917 3644 1923
rect 3796 1917 3820 1923
rect 3860 1917 3980 1923
rect 4148 1917 4163 1923
rect 4045 1904 4051 1916
rect 3453 1897 3516 1903
rect 3540 1897 3564 1903
rect 3604 1897 4035 1903
rect 180 1877 364 1883
rect 372 1877 796 1883
rect 852 1877 972 1883
rect 1012 1877 1068 1883
rect 1108 1877 1132 1883
rect 1300 1877 1308 1883
rect 1332 1877 1468 1883
rect 1501 1877 1644 1883
rect 180 1857 220 1863
rect 772 1857 876 1863
rect 884 1857 1100 1863
rect 1236 1857 1283 1863
rect 196 1837 252 1843
rect 260 1837 396 1843
rect 596 1837 620 1843
rect 644 1837 668 1843
rect 852 1837 1260 1843
rect 1277 1843 1283 1857
rect 1325 1863 1331 1876
rect 1501 1863 1507 1877
rect 1652 1877 1708 1883
rect 1780 1877 2092 1883
rect 2164 1877 2268 1883
rect 2292 1877 2316 1883
rect 2340 1877 2348 1883
rect 2372 1877 2403 1883
rect 1300 1857 1331 1863
rect 1453 1857 1507 1863
rect 1277 1837 1420 1843
rect 564 1817 652 1823
rect 660 1817 684 1823
rect 708 1817 1068 1823
rect 1092 1817 1132 1823
rect 1172 1817 1228 1823
rect 1252 1817 1292 1823
rect 1332 1817 1340 1823
rect 1453 1823 1459 1857
rect 1556 1857 1676 1863
rect 1684 1857 1836 1863
rect 1853 1857 1884 1863
rect 1652 1837 1667 1843
rect 1444 1817 1459 1823
rect 1476 1817 1548 1823
rect 1661 1823 1667 1837
rect 1684 1837 1772 1843
rect 1853 1843 1859 1857
rect 1924 1857 1980 1863
rect 2004 1857 2204 1863
rect 2260 1857 2380 1863
rect 2397 1863 2403 1877
rect 2436 1877 2460 1883
rect 2484 1877 2636 1883
rect 2740 1877 2764 1883
rect 2772 1877 2812 1883
rect 2900 1877 2956 1883
rect 3060 1877 3260 1883
rect 3284 1877 3340 1883
rect 3348 1877 3388 1883
rect 3412 1877 3548 1883
rect 3572 1877 3804 1883
rect 3828 1877 3884 1883
rect 3988 1877 4012 1883
rect 4029 1883 4035 1897
rect 4116 1897 4140 1903
rect 4157 1903 4163 1917
rect 4244 1917 4332 1923
rect 4340 1917 4572 1923
rect 4612 1917 4844 1923
rect 4916 1917 4924 1923
rect 4932 1917 4940 1923
rect 5108 1917 5548 1923
rect 5556 1917 5580 1923
rect 5668 1917 5820 1923
rect 5988 1917 6060 1923
rect 6116 1917 6252 1923
rect 5069 1904 5075 1916
rect 4157 1897 4172 1903
rect 4196 1897 4204 1903
rect 4212 1897 4268 1903
rect 4388 1897 4460 1903
rect 4532 1897 4540 1903
rect 4612 1897 4620 1903
rect 4660 1897 4748 1903
rect 4772 1897 4828 1903
rect 4868 1897 4876 1903
rect 5300 1897 5372 1903
rect 5380 1897 5436 1903
rect 5716 1897 5996 1903
rect 6036 1897 6140 1903
rect 6212 1897 6252 1903
rect 6253 1884 6259 1896
rect 4029 1877 4060 1883
rect 4212 1877 4332 1883
rect 4340 1877 4444 1883
rect 4452 1877 5084 1883
rect 5092 1877 5148 1883
rect 5316 1877 5324 1883
rect 5396 1877 5452 1883
rect 5684 1877 5772 1883
rect 6084 1877 6124 1883
rect 6180 1877 6236 1883
rect 2397 1857 2627 1863
rect 1796 1837 1859 1843
rect 1956 1837 1980 1843
rect 2004 1837 2035 1843
rect 1661 1817 1692 1823
rect 1716 1817 1740 1823
rect 1796 1817 1820 1823
rect 1860 1817 2012 1823
rect 2029 1823 2035 1837
rect 2052 1837 2076 1843
rect 2100 1837 2284 1843
rect 2301 1837 2380 1843
rect 2029 1817 2140 1823
rect 2164 1817 2172 1823
rect 2301 1823 2307 1837
rect 2420 1837 2540 1843
rect 2564 1837 2604 1843
rect 2621 1843 2627 1857
rect 2788 1857 2812 1863
rect 3220 1857 3267 1863
rect 2621 1837 2691 1843
rect 2196 1817 2307 1823
rect 2388 1817 2444 1823
rect 2580 1817 2668 1823
rect 2685 1823 2691 1837
rect 2740 1837 2764 1843
rect 2820 1837 2972 1843
rect 3028 1837 3212 1843
rect 3261 1843 3267 1857
rect 3284 1857 3308 1863
rect 3348 1857 3372 1863
rect 3380 1857 3596 1863
rect 3668 1857 3724 1863
rect 3748 1857 4124 1863
rect 4148 1857 4380 1863
rect 4436 1857 4803 1863
rect 3261 1837 3308 1843
rect 3380 1837 3491 1843
rect 2685 1817 2732 1823
rect 3268 1817 3276 1823
rect 3300 1817 3324 1823
rect 3380 1817 3468 1823
rect 3485 1823 3491 1837
rect 3636 1837 3692 1843
rect 3700 1837 4028 1843
rect 4036 1837 4556 1843
rect 4564 1837 4620 1843
rect 4628 1837 4764 1843
rect 4772 1837 4780 1843
rect 4797 1843 4803 1857
rect 4852 1857 4860 1863
rect 4868 1857 5100 1863
rect 5140 1857 5260 1863
rect 5460 1857 5500 1863
rect 5716 1857 5724 1863
rect 5940 1857 6028 1863
rect 6196 1857 6268 1863
rect 4797 1837 5724 1843
rect 5908 1837 5964 1843
rect 5972 1837 6012 1843
rect 3485 1817 3852 1823
rect 3908 1817 4044 1823
rect 4100 1817 4140 1823
rect 4189 1817 4572 1823
rect 3112 1814 3160 1816
rect 484 1797 620 1803
rect 644 1797 716 1803
rect 724 1797 1196 1803
rect 1220 1797 1276 1803
rect 1380 1797 1420 1803
rect 1460 1797 1484 1803
rect 1508 1797 1619 1803
rect 436 1777 604 1783
rect 612 1777 860 1783
rect 1044 1777 1068 1783
rect 1108 1777 1292 1783
rect 1613 1783 1619 1797
rect 1636 1797 1660 1803
rect 1741 1797 2028 1803
rect 1741 1783 1747 1797
rect 2036 1797 2044 1803
rect 2132 1797 2156 1803
rect 2196 1797 2348 1803
rect 2372 1797 2460 1803
rect 2548 1797 2572 1803
rect 2596 1797 2876 1803
rect 3112 1806 3113 1814
rect 3122 1806 3123 1814
rect 3158 1806 3160 1814
rect 3112 1804 3160 1806
rect 2964 1800 3020 1803
rect 2957 1797 3020 1800
rect 3220 1797 3292 1803
rect 3332 1797 3356 1803
rect 3396 1797 3420 1803
rect 3444 1797 3532 1803
rect 3540 1797 3660 1803
rect 3700 1797 3724 1803
rect 3764 1797 3836 1803
rect 4189 1803 4195 1817
rect 4820 1817 4844 1823
rect 4900 1817 4908 1823
rect 5124 1817 5244 1823
rect 5252 1817 5484 1823
rect 5508 1817 5612 1823
rect 6020 1817 6028 1823
rect 6116 1817 6204 1823
rect 3860 1797 4195 1803
rect 4212 1797 4236 1803
rect 4292 1797 4316 1803
rect 4340 1797 4524 1803
rect 4596 1797 4652 1803
rect 4724 1797 5868 1803
rect 5988 1797 6220 1803
rect 1613 1777 1747 1783
rect 1876 1777 2060 1783
rect 2084 1777 2252 1783
rect 2292 1777 2380 1783
rect 2484 1780 2700 1783
rect 2477 1777 2700 1780
rect 2724 1777 2796 1783
rect 2852 1780 2963 1783
rect 2852 1777 2956 1780
rect 2973 1777 3084 1783
rect 2973 1764 2979 1777
rect 3204 1777 3580 1783
rect 3588 1777 4220 1783
rect 4228 1777 4700 1783
rect 4884 1777 4988 1783
rect 5012 1777 5052 1783
rect 5444 1777 5516 1783
rect 5524 1777 5532 1783
rect 5620 1777 5644 1783
rect 5796 1777 6188 1783
rect 68 1757 76 1763
rect 244 1757 332 1763
rect 340 1757 476 1763
rect 484 1757 508 1763
rect 676 1757 716 1763
rect 724 1757 828 1763
rect 948 1757 1100 1763
rect 1524 1757 1811 1763
rect 36 1737 124 1743
rect 132 1737 172 1743
rect 468 1737 764 1743
rect 820 1737 1052 1743
rect 1172 1737 1244 1743
rect 1252 1737 1740 1743
rect 1805 1743 1811 1757
rect 1940 1757 1996 1763
rect 2052 1757 2156 1763
rect 2164 1757 2348 1763
rect 2397 1760 2483 1763
rect 2397 1757 2476 1760
rect 1805 1737 1852 1743
rect 1908 1737 1948 1743
rect 2036 1737 2060 1743
rect 2132 1737 2156 1743
rect 2212 1737 2300 1743
rect 2324 1737 2339 1743
rect 20 1717 108 1723
rect 324 1717 492 1723
rect 596 1717 620 1723
rect 692 1717 748 1723
rect 820 1717 860 1723
rect 1028 1717 1324 1723
rect 1380 1717 1420 1723
rect 1492 1717 1708 1723
rect 1716 1717 1836 1723
rect 1892 1717 1900 1723
rect 1956 1717 1964 1723
rect 1988 1717 2220 1723
rect 2244 1717 2284 1723
rect 2292 1717 2316 1723
rect 2333 1723 2339 1737
rect 2397 1743 2403 1757
rect 2548 1757 2588 1763
rect 2772 1757 2972 1763
rect 2996 1757 3084 1763
rect 3364 1757 3388 1763
rect 3428 1757 3500 1763
rect 3572 1757 3612 1763
rect 3620 1757 3676 1763
rect 3684 1757 3692 1763
rect 3732 1757 3772 1763
rect 3796 1757 3804 1763
rect 3812 1757 3900 1763
rect 3988 1757 3996 1763
rect 4020 1757 4364 1763
rect 4420 1757 5468 1763
rect 5476 1757 5516 1763
rect 5540 1757 5580 1763
rect 5604 1757 5724 1763
rect 5876 1757 6076 1763
rect 2356 1737 2403 1743
rect 2420 1737 2508 1743
rect 2708 1737 2796 1743
rect 2836 1737 2860 1743
rect 2948 1737 2956 1743
rect 2996 1737 3500 1743
rect 3508 1737 3932 1743
rect 3940 1737 4268 1743
rect 4324 1737 4332 1743
rect 4564 1737 4684 1743
rect 5044 1737 5068 1743
rect 5076 1737 5084 1743
rect 5268 1737 5324 1743
rect 5476 1737 5820 1743
rect 5828 1737 5836 1743
rect 2333 1717 2412 1723
rect 2436 1717 2444 1723
rect 2452 1717 2556 1723
rect 2564 1717 2876 1723
rect 3396 1717 3468 1723
rect 3508 1717 3740 1723
rect 3764 1717 3820 1723
rect 4276 1717 5612 1723
rect 5636 1717 5692 1723
rect 5732 1717 5836 1723
rect 6036 1717 6140 1723
rect 1325 1704 1331 1716
rect 116 1697 156 1703
rect 180 1697 204 1703
rect 436 1697 588 1703
rect 1076 1697 1196 1703
rect 1348 1697 1372 1703
rect 1437 1697 1516 1703
rect 468 1677 732 1683
rect 1437 1683 1443 1697
rect 1812 1697 1868 1703
rect 1924 1697 2012 1703
rect 2100 1697 2124 1703
rect 2164 1697 2700 1703
rect 2724 1697 2780 1703
rect 2804 1697 2860 1703
rect 2900 1697 3820 1703
rect 3940 1697 3964 1703
rect 3997 1697 4108 1703
rect 788 1677 1443 1683
rect 1476 1677 1516 1683
rect 1556 1677 1964 1683
rect 2004 1677 2092 1683
rect 2228 1677 2380 1683
rect 2452 1677 2540 1683
rect 2557 1677 2604 1683
rect 724 1657 796 1663
rect 836 1657 892 1663
rect 916 1657 1027 1663
rect 308 1637 1004 1643
rect 1021 1643 1027 1657
rect 1044 1657 1132 1663
rect 1140 1657 1260 1663
rect 1396 1657 1740 1663
rect 1892 1657 1932 1663
rect 1972 1657 2060 1663
rect 2116 1657 2204 1663
rect 2228 1657 2396 1663
rect 2557 1663 2563 1677
rect 2628 1677 2636 1683
rect 2772 1677 2812 1683
rect 2836 1677 2844 1683
rect 2932 1677 3212 1683
rect 3236 1677 3244 1683
rect 3997 1683 4003 1697
rect 4180 1697 4188 1703
rect 4308 1697 4428 1703
rect 4452 1697 4476 1703
rect 4500 1697 4716 1703
rect 4804 1697 5196 1703
rect 5204 1697 5276 1703
rect 5300 1697 5388 1703
rect 5460 1697 5532 1703
rect 5620 1697 5660 1703
rect 5988 1697 6252 1703
rect 3268 1677 4003 1683
rect 4020 1677 4108 1683
rect 4132 1677 4220 1683
rect 4237 1677 4924 1683
rect 2420 1657 2563 1663
rect 2756 1657 2892 1663
rect 4237 1663 4243 1677
rect 5444 1677 5596 1683
rect 2916 1657 4243 1663
rect 4260 1657 4300 1663
rect 4388 1657 4652 1663
rect 4756 1657 4812 1663
rect 4916 1657 5148 1663
rect 5588 1657 5612 1663
rect 5812 1657 5836 1663
rect 1021 1637 1052 1643
rect 1076 1637 1996 1643
rect 2004 1637 2540 1643
rect 2548 1637 3404 1643
rect 3412 1637 4860 1643
rect 4868 1637 5004 1643
rect 5012 1637 5036 1643
rect 5076 1637 5484 1643
rect 5572 1637 5596 1643
rect 5876 1637 5884 1643
rect 5892 1637 5964 1643
rect 532 1617 876 1623
rect 964 1617 1068 1623
rect 1108 1617 1148 1623
rect 1156 1617 1244 1623
rect 1268 1617 1276 1623
rect 1364 1617 1532 1623
rect 1652 1617 2588 1623
rect 2612 1617 2668 1623
rect 2692 1617 2716 1623
rect 2804 1617 2828 1623
rect 2868 1617 2892 1623
rect 2932 1617 4012 1623
rect 4148 1617 4252 1623
rect 4276 1617 4572 1623
rect 4596 1617 4643 1623
rect 1576 1614 1624 1616
rect 1576 1606 1577 1614
rect 1586 1606 1587 1614
rect 1622 1606 1624 1614
rect 1576 1604 1624 1606
rect 4637 1604 4643 1617
rect 4852 1617 4956 1623
rect 5092 1617 5276 1623
rect 5396 1617 6140 1623
rect 4664 1614 4712 1616
rect 4664 1606 4665 1614
rect 4674 1606 4675 1614
rect 4710 1606 4712 1614
rect 4664 1604 4712 1606
rect 980 1597 1244 1603
rect 1332 1597 1379 1603
rect 676 1577 748 1583
rect 756 1577 764 1583
rect 1012 1577 1356 1583
rect 1373 1583 1379 1597
rect 1476 1597 1516 1603
rect 1652 1597 1708 1603
rect 1764 1597 1916 1603
rect 1940 1597 2044 1603
rect 2100 1597 2220 1603
rect 2308 1597 2348 1603
rect 2372 1597 2572 1603
rect 2596 1597 2860 1603
rect 2868 1597 2924 1603
rect 3588 1597 3612 1603
rect 3636 1597 3756 1603
rect 3924 1597 4236 1603
rect 4308 1597 4460 1603
rect 4500 1597 4588 1603
rect 4740 1597 5836 1603
rect 6164 1597 6268 1603
rect 1373 1577 1660 1583
rect 1700 1577 1868 1583
rect 1972 1577 1980 1583
rect 1988 1577 2028 1583
rect 2100 1577 2156 1583
rect 2180 1577 3452 1583
rect 3476 1577 3548 1583
rect 3572 1577 4012 1583
rect 4212 1577 4332 1583
rect 4372 1577 4492 1583
rect 4580 1577 4668 1583
rect 4692 1577 5468 1583
rect 5492 1577 5660 1583
rect 5812 1577 5980 1583
rect 324 1557 492 1563
rect 788 1557 812 1563
rect 884 1557 1036 1563
rect 1181 1557 2451 1563
rect 276 1537 364 1543
rect 548 1537 940 1543
rect 996 1537 1100 1543
rect 1181 1543 1187 1557
rect 1140 1537 1187 1543
rect 1236 1537 1292 1543
rect 1332 1537 1548 1543
rect 1661 1537 1740 1543
rect -19 1517 300 1523
rect 404 1517 428 1523
rect 580 1517 732 1523
rect 756 1517 771 1523
rect 52 1497 220 1503
rect 228 1497 236 1503
rect 253 1497 428 1503
rect 253 1483 259 1497
rect 564 1497 700 1503
rect 724 1497 748 1503
rect 212 1477 259 1483
rect 276 1477 332 1483
rect 340 1477 364 1483
rect 765 1483 771 1517
rect 820 1517 844 1523
rect 852 1517 940 1523
rect 973 1517 1052 1523
rect 788 1497 867 1503
rect 765 1477 796 1483
rect 861 1483 867 1497
rect 973 1503 979 1517
rect 1060 1517 1084 1523
rect 1140 1517 1196 1523
rect 1236 1517 1260 1523
rect 1300 1517 1404 1523
rect 1428 1517 1468 1523
rect 1492 1517 1500 1523
rect 1661 1523 1667 1537
rect 1764 1537 1804 1543
rect 1844 1537 2124 1543
rect 2148 1537 2268 1543
rect 2292 1537 2380 1543
rect 2445 1543 2451 1557
rect 2484 1557 2499 1563
rect 2445 1537 2476 1543
rect 2493 1543 2499 1557
rect 2564 1557 2588 1563
rect 2605 1557 2652 1563
rect 2605 1543 2611 1557
rect 2708 1557 3468 1563
rect 3668 1557 3724 1563
rect 3796 1557 3900 1563
rect 3924 1557 4204 1563
rect 4324 1557 4556 1563
rect 4596 1557 5043 1563
rect 2493 1537 2611 1543
rect 2644 1537 2732 1543
rect 2772 1537 3100 1543
rect 3124 1537 3244 1543
rect 3268 1537 3436 1543
rect 3444 1537 3500 1543
rect 3572 1537 4252 1543
rect 4276 1537 4364 1543
rect 4404 1537 4428 1543
rect 4468 1537 4851 1543
rect 1540 1517 1667 1523
rect 1684 1517 1820 1523
rect 1940 1517 1964 1523
rect 2020 1517 2092 1523
rect 2116 1517 2140 1523
rect 2244 1517 2316 1523
rect 2340 1517 2396 1523
rect 2420 1517 2764 1523
rect 2804 1517 2844 1523
rect 2980 1517 3020 1523
rect 3092 1517 3132 1523
rect 3316 1517 3932 1523
rect 3988 1517 4323 1523
rect 884 1497 979 1503
rect 996 1497 1020 1503
rect 1028 1497 1052 1503
rect 1108 1497 1244 1503
rect 1268 1497 1395 1503
rect 861 1477 876 1483
rect 900 1477 1132 1483
rect 1156 1477 1212 1483
rect 1236 1477 1260 1483
rect 1389 1483 1395 1497
rect 1428 1497 1452 1503
rect 1476 1497 1587 1503
rect 1389 1477 1436 1483
rect 1581 1483 1587 1497
rect 1604 1497 1644 1503
rect 1652 1497 1676 1503
rect 1748 1497 2044 1503
rect 2068 1497 2268 1503
rect 2308 1497 2364 1503
rect 2388 1497 2460 1503
rect 2468 1497 2492 1503
rect 2516 1497 2780 1503
rect 2820 1497 2963 1503
rect 1453 1477 1507 1483
rect 1581 1477 1772 1483
rect 420 1457 812 1463
rect 580 1437 604 1443
rect 708 1437 780 1443
rect 829 1443 835 1476
rect 852 1457 988 1463
rect 1012 1457 1196 1463
rect 1268 1457 1388 1463
rect 1396 1457 1420 1463
rect 1453 1463 1459 1477
rect 1428 1457 1459 1463
rect 1501 1463 1507 1477
rect 1876 1477 2028 1483
rect 2068 1477 2092 1483
rect 2132 1477 2188 1483
rect 2292 1477 2348 1483
rect 2484 1477 2643 1483
rect 1501 1457 1532 1463
rect 1540 1457 1596 1463
rect 1668 1457 1724 1463
rect 1780 1457 1900 1463
rect 1924 1457 1948 1463
rect 2052 1457 2140 1463
rect 2164 1457 2188 1463
rect 2436 1457 2492 1463
rect 2516 1457 2524 1463
rect 2580 1457 2588 1463
rect 2637 1463 2643 1477
rect 2660 1477 2700 1483
rect 2797 1483 2803 1496
rect 2724 1477 2803 1483
rect 2836 1477 2892 1483
rect 2932 1477 2940 1483
rect 2957 1483 2963 1497
rect 3108 1497 3372 1503
rect 3572 1497 3628 1503
rect 3716 1497 3916 1503
rect 3956 1497 4012 1503
rect 4132 1497 4300 1503
rect 4317 1503 4323 1517
rect 4404 1517 4732 1523
rect 4772 1517 4828 1523
rect 4845 1523 4851 1537
rect 4868 1537 5020 1543
rect 5037 1543 5043 1557
rect 5172 1557 5260 1563
rect 5268 1557 5756 1563
rect 5780 1557 5820 1563
rect 5844 1557 6108 1563
rect 5037 1537 5196 1543
rect 5268 1537 5948 1543
rect 6020 1537 6220 1543
rect 6237 1537 6252 1543
rect 4845 1517 4876 1523
rect 4884 1517 4956 1523
rect 5220 1517 5292 1523
rect 5316 1517 5340 1523
rect 5508 1517 5548 1523
rect 5764 1517 5772 1523
rect 5956 1517 6044 1523
rect 6237 1523 6243 1537
rect 6189 1517 6243 1523
rect 4317 1500 4460 1503
rect 4317 1497 4467 1500
rect 5028 1497 5068 1503
rect 5252 1497 5516 1503
rect 5524 1497 5532 1503
rect 5588 1497 5676 1503
rect 5716 1497 5740 1503
rect 5748 1497 5804 1503
rect 5812 1497 5932 1503
rect 5956 1497 6012 1503
rect 6068 1497 6076 1503
rect 4813 1484 4819 1496
rect 4941 1484 4947 1496
rect 2957 1477 3196 1483
rect 3220 1477 3260 1483
rect 3316 1477 3404 1483
rect 3460 1477 3468 1483
rect 3565 1477 3644 1483
rect 3565 1464 3571 1477
rect 3860 1477 3932 1483
rect 4052 1477 4268 1483
rect 4292 1477 4348 1483
rect 4461 1480 4524 1483
rect 4468 1477 4524 1480
rect 4596 1477 4611 1483
rect 2637 1457 2764 1463
rect 2804 1457 2988 1463
rect 3012 1457 3036 1463
rect 3108 1457 3164 1463
rect 3236 1457 3340 1463
rect 3380 1457 3452 1463
rect 3460 1457 3532 1463
rect 3636 1457 4396 1463
rect 4468 1457 4588 1463
rect 4605 1463 4611 1477
rect 4644 1477 4748 1483
rect 4836 1477 4908 1483
rect 5044 1477 5260 1483
rect 5332 1477 5404 1483
rect 5428 1477 5548 1483
rect 5780 1477 5836 1483
rect 5860 1477 5996 1483
rect 6004 1477 6028 1483
rect 6036 1477 6092 1483
rect 6189 1483 6195 1517
rect 6212 1497 6252 1503
rect 6180 1477 6195 1483
rect 4605 1457 4668 1463
rect 4701 1457 5132 1463
rect 813 1437 835 1443
rect 324 1417 748 1423
rect 756 1417 764 1423
rect 813 1423 819 1437
rect 868 1437 1228 1443
rect 1268 1437 1340 1443
rect 1348 1437 1676 1443
rect 1780 1437 1900 1443
rect 1956 1437 2060 1443
rect 2189 1437 2892 1443
rect 788 1417 819 1423
rect 836 1417 844 1423
rect 852 1417 860 1423
rect 884 1417 1004 1423
rect 1012 1417 1020 1423
rect 1044 1417 1116 1423
rect 1172 1417 1228 1423
rect 1364 1417 1404 1423
rect 1412 1417 1516 1423
rect 1604 1417 1740 1423
rect 2189 1423 2195 1437
rect 2948 1437 3020 1443
rect 3204 1437 3308 1443
rect 3444 1437 3468 1443
rect 3524 1437 3788 1443
rect 3812 1437 4188 1443
rect 4212 1437 4412 1443
rect 4701 1443 4707 1457
rect 5252 1457 5292 1463
rect 5332 1457 5420 1463
rect 5428 1457 5580 1463
rect 5588 1457 5724 1463
rect 5732 1457 5788 1463
rect 5796 1457 5836 1463
rect 5844 1457 5916 1463
rect 6100 1457 6124 1463
rect 4564 1437 4707 1443
rect 4724 1437 4860 1443
rect 4884 1437 5484 1443
rect 5652 1437 5932 1443
rect 1812 1417 2195 1423
rect 2260 1417 2332 1423
rect 2356 1417 2428 1423
rect 2612 1417 2668 1423
rect 2708 1417 2764 1423
rect 2772 1417 2876 1423
rect 2884 1417 3004 1423
rect 3220 1417 3388 1423
rect 3412 1417 3660 1423
rect 4052 1417 4140 1423
rect 4164 1417 4892 1423
rect 4900 1417 5052 1423
rect 5060 1417 5100 1423
rect 5108 1417 5308 1423
rect 5316 1417 5452 1423
rect 5684 1417 5916 1423
rect 5972 1417 6028 1423
rect 6036 1417 6204 1423
rect 3112 1414 3160 1416
rect 3112 1406 3113 1414
rect 3122 1406 3123 1414
rect 3158 1406 3160 1414
rect 3112 1404 3160 1406
rect 612 1397 908 1403
rect 1060 1397 1100 1403
rect 1140 1397 1612 1403
rect 1636 1397 1676 1403
rect 1748 1397 1836 1403
rect 1892 1397 2028 1403
rect 2100 1397 2172 1403
rect 2196 1397 2364 1403
rect 2381 1397 2828 1403
rect 68 1377 236 1383
rect 244 1377 844 1383
rect 852 1377 940 1383
rect 948 1377 956 1383
rect 980 1377 1228 1383
rect 1300 1377 1580 1383
rect 2381 1383 2387 1397
rect 2836 1397 3068 1403
rect 3188 1397 3292 1403
rect 3380 1397 3436 1403
rect 3460 1397 3900 1403
rect 3924 1397 3932 1403
rect 3940 1397 4076 1403
rect 4148 1397 4172 1403
rect 4244 1397 4252 1403
rect 4276 1397 4556 1403
rect 4660 1397 4780 1403
rect 4836 1397 4844 1403
rect 4996 1397 5772 1403
rect 5780 1397 5804 1403
rect 5940 1397 5964 1403
rect 4109 1384 4115 1396
rect 1620 1377 2387 1383
rect 2404 1377 2636 1383
rect 2644 1377 2780 1383
rect 2788 1377 2860 1383
rect 2916 1377 2972 1383
rect 2996 1377 3011 1383
rect 164 1357 332 1363
rect 340 1357 476 1363
rect 484 1357 652 1363
rect 660 1357 748 1363
rect 772 1357 899 1363
rect 196 1337 268 1343
rect 308 1337 316 1343
rect 420 1337 508 1343
rect 532 1337 588 1343
rect 628 1337 876 1343
rect 893 1343 899 1357
rect 948 1357 1356 1363
rect 1396 1357 1404 1363
rect 1428 1357 1436 1363
rect 1460 1357 1484 1363
rect 1556 1357 1612 1363
rect 1668 1357 1804 1363
rect 1844 1357 1852 1363
rect 1876 1357 1900 1363
rect 2036 1357 2108 1363
rect 2196 1357 2252 1363
rect 2308 1357 2316 1363
rect 2388 1357 2652 1363
rect 2660 1357 2828 1363
rect 2836 1357 2988 1363
rect 3005 1363 3011 1377
rect 3028 1377 3132 1383
rect 3156 1377 3212 1383
rect 3428 1377 3532 1383
rect 3764 1377 3980 1383
rect 4228 1377 4316 1383
rect 4340 1377 4492 1383
rect 4580 1377 4668 1383
rect 4676 1377 4844 1383
rect 4868 1377 4924 1383
rect 5060 1377 5628 1383
rect 5844 1377 5996 1383
rect 6084 1377 6188 1383
rect 3629 1364 3635 1376
rect 3005 1357 3084 1363
rect 3124 1357 3523 1363
rect 893 1337 1020 1343
rect 1044 1337 1084 1343
rect 1108 1337 1164 1343
rect 1268 1337 1372 1343
rect 1396 1337 1436 1343
rect 1492 1337 1548 1343
rect 1572 1337 1612 1343
rect 1652 1337 1788 1343
rect 2036 1337 2211 1343
rect -19 1317 12 1323
rect 180 1317 220 1323
rect 269 1323 275 1336
rect 269 1317 444 1323
rect 724 1317 796 1323
rect 804 1317 876 1323
rect 900 1317 956 1323
rect 964 1317 1164 1323
rect 1220 1317 1292 1323
rect 1300 1317 1484 1323
rect 1540 1317 1660 1323
rect 1748 1317 1820 1323
rect 1892 1317 1964 1323
rect 2020 1317 2076 1323
rect 2164 1317 2188 1323
rect 2205 1323 2211 1337
rect 2228 1337 2316 1343
rect 2356 1337 2483 1343
rect 2205 1317 2380 1323
rect 2436 1317 2444 1323
rect 2477 1323 2483 1337
rect 2500 1337 2652 1343
rect 2676 1337 2684 1343
rect 2708 1337 2796 1343
rect 2804 1337 2812 1343
rect 2829 1337 2844 1343
rect 2477 1317 2556 1323
rect 2580 1317 2620 1323
rect 2644 1317 2700 1323
rect 2724 1317 2764 1323
rect 2829 1323 2835 1337
rect 2852 1337 3020 1343
rect 3172 1337 3372 1343
rect 3396 1337 3436 1343
rect 3517 1343 3523 1357
rect 3668 1357 3676 1363
rect 4084 1357 4092 1363
rect 4100 1357 4172 1363
rect 4404 1357 4956 1363
rect 4964 1357 5004 1363
rect 5060 1357 5196 1363
rect 5348 1357 5836 1363
rect 5908 1357 6028 1363
rect 3517 1337 3788 1343
rect 3892 1337 4012 1343
rect 4100 1337 4108 1343
rect 4148 1337 4348 1343
rect 4516 1337 4652 1343
rect 4756 1337 4988 1343
rect 4996 1337 5020 1343
rect 5044 1337 5276 1343
rect 5540 1337 5676 1343
rect 5716 1337 5964 1343
rect 6004 1337 6044 1343
rect 2788 1317 2835 1323
rect 2852 1317 2876 1323
rect 2980 1317 2988 1323
rect 3252 1317 3276 1323
rect 3300 1317 3500 1323
rect 3540 1317 3692 1323
rect 3812 1317 3980 1323
rect 4068 1317 4220 1323
rect 4276 1317 4844 1323
rect 4852 1317 5132 1323
rect 5236 1317 5308 1323
rect 5364 1317 5372 1323
rect 5524 1317 5532 1323
rect 5581 1317 5612 1323
rect 3181 1304 3187 1316
rect 772 1297 892 1303
rect 932 1297 1004 1303
rect 1092 1297 1116 1303
rect 1156 1297 1212 1303
rect 1252 1297 1356 1303
rect 1380 1297 1436 1303
rect 1508 1297 1596 1303
rect 1620 1297 1708 1303
rect 1773 1297 2028 1303
rect 372 1277 1164 1283
rect 1220 1277 1260 1283
rect 1332 1277 1404 1283
rect 1444 1277 1532 1283
rect 1773 1283 1779 1297
rect 2068 1297 2172 1303
rect 2180 1297 2412 1303
rect 2500 1297 2524 1303
rect 2532 1297 2588 1303
rect 2612 1297 3052 1303
rect 3284 1297 3340 1303
rect 3380 1297 3420 1303
rect 3476 1297 3916 1303
rect 4020 1297 4316 1303
rect 4404 1297 4476 1303
rect 4532 1297 4540 1303
rect 4772 1297 4860 1303
rect 4900 1297 4924 1303
rect 4948 1297 5004 1303
rect 5028 1297 5132 1303
rect 1549 1277 1779 1283
rect 708 1257 1036 1263
rect 1060 1257 1196 1263
rect 1316 1257 1356 1263
rect 1549 1263 1555 1277
rect 1844 1277 1948 1283
rect 1972 1277 2060 1283
rect 2132 1277 2348 1283
rect 2388 1277 2508 1283
rect 2596 1277 2620 1283
rect 2644 1277 2652 1283
rect 2788 1277 2796 1283
rect 2820 1277 2828 1283
rect 2868 1277 2892 1283
rect 2900 1277 3020 1283
rect 3044 1277 3164 1283
rect 3188 1277 3372 1283
rect 3492 1277 3500 1283
rect 3540 1277 3660 1283
rect 3860 1277 4316 1283
rect 4324 1277 4556 1283
rect 4596 1277 4716 1283
rect 4788 1277 4876 1283
rect 4916 1277 5212 1283
rect 5316 1277 5452 1283
rect 5581 1264 5587 1317
rect 5812 1317 6012 1323
rect 6068 1317 6108 1323
rect 5597 1297 5724 1303
rect 1492 1257 1555 1263
rect 1652 1257 1852 1263
rect 1924 1257 2028 1263
rect 2100 1257 2444 1263
rect 2452 1257 3244 1263
rect 3252 1257 3276 1263
rect 3300 1257 3388 1263
rect 3412 1257 3596 1263
rect 4340 1257 5020 1263
rect 5076 1257 5404 1263
rect 308 1237 716 1243
rect 724 1237 1100 1243
rect 1108 1237 1132 1243
rect 1188 1237 1324 1243
rect 1364 1237 1436 1243
rect 1460 1237 1900 1243
rect 2045 1237 2108 1243
rect 164 1217 556 1223
rect 564 1217 812 1223
rect 820 1217 1004 1223
rect 1012 1217 1036 1223
rect 1124 1217 1468 1223
rect 1524 1217 1548 1223
rect 2045 1223 2051 1237
rect 2132 1237 2268 1243
rect 2292 1237 2348 1243
rect 2372 1237 2412 1243
rect 2452 1237 2588 1243
rect 2612 1237 3596 1243
rect 3684 1237 3820 1243
rect 3828 1237 3964 1243
rect 3972 1237 4028 1243
rect 4036 1237 4252 1243
rect 4260 1237 4300 1243
rect 4308 1237 4348 1243
rect 4420 1237 4492 1243
rect 4516 1237 4972 1243
rect 5092 1237 5100 1243
rect 5300 1237 5340 1243
rect 5597 1243 5603 1297
rect 5757 1297 5916 1303
rect 5757 1283 5763 1297
rect 6036 1297 6188 1303
rect 5732 1277 5763 1283
rect 5908 1277 5980 1283
rect 6068 1277 6140 1283
rect 6196 1277 6268 1283
rect 5700 1257 6268 1263
rect 5588 1237 5603 1243
rect 5956 1237 5996 1243
rect 1684 1217 2051 1223
rect 2068 1217 2220 1223
rect 2260 1217 2307 1223
rect 740 1197 924 1203
rect 1012 1197 1260 1203
rect 1300 1197 1404 1203
rect 1469 1203 1475 1216
rect 1576 1214 1624 1216
rect 1576 1206 1577 1214
rect 1586 1206 1587 1214
rect 1622 1206 1624 1214
rect 1576 1204 1624 1206
rect 1469 1197 1548 1203
rect 1709 1197 1804 1203
rect 84 1177 124 1183
rect 132 1177 284 1183
rect 580 1177 716 1183
rect 932 1177 940 1183
rect 1076 1177 1132 1183
rect 1709 1183 1715 1197
rect 1876 1197 2220 1203
rect 2260 1197 2284 1203
rect 2301 1203 2307 1217
rect 2324 1217 2364 1223
rect 2484 1217 2540 1223
rect 2564 1217 2940 1223
rect 2980 1217 3564 1223
rect 3732 1217 4380 1223
rect 4500 1217 4588 1223
rect 4788 1217 5068 1223
rect 5156 1217 5164 1223
rect 5220 1217 5308 1223
rect 5492 1217 5612 1223
rect 5828 1217 6060 1223
rect 4664 1214 4712 1216
rect 4664 1206 4665 1214
rect 4674 1206 4675 1214
rect 4710 1206 4712 1214
rect 4664 1204 4712 1206
rect 2301 1197 2380 1203
rect 2436 1197 2732 1203
rect 2749 1197 2796 1203
rect 1172 1177 1715 1183
rect 1732 1177 1804 1183
rect 2052 1177 2156 1183
rect 2180 1177 2300 1183
rect 2324 1177 2700 1183
rect 2749 1183 2755 1197
rect 2820 1197 3148 1203
rect 3172 1197 3212 1203
rect 3572 1197 3724 1203
rect 3924 1197 4092 1203
rect 4100 1197 4556 1203
rect 4756 1197 5331 1203
rect 2740 1177 2755 1183
rect 2804 1177 3084 1183
rect 3140 1177 3196 1183
rect 3220 1177 3756 1183
rect 4340 1177 4508 1183
rect 4532 1177 4732 1183
rect 4836 1177 5180 1183
rect 5325 1183 5331 1197
rect 5524 1197 5596 1203
rect 5780 1197 5868 1203
rect 5940 1197 6012 1203
rect 6141 1197 6188 1203
rect 5325 1177 5676 1183
rect 5876 1177 5900 1183
rect 6141 1183 6147 1197
rect 6212 1197 6220 1203
rect 5972 1177 6147 1183
rect 6180 1177 6220 1183
rect 292 1157 412 1163
rect 676 1157 684 1163
rect 692 1157 732 1163
rect 756 1157 2636 1163
rect 2660 1157 2700 1163
rect 2724 1157 3052 1163
rect 3076 1157 3612 1163
rect 3620 1157 3836 1163
rect 3892 1157 4108 1163
rect 4116 1157 4284 1163
rect 4308 1157 4412 1163
rect 4436 1157 4668 1163
rect 5140 1157 5260 1163
rect 5268 1157 5340 1163
rect 5348 1157 5564 1163
rect 5572 1157 5676 1163
rect 5844 1157 6220 1163
rect 500 1137 588 1143
rect 596 1137 700 1143
rect 724 1137 748 1143
rect 772 1137 812 1143
rect 1060 1137 1244 1143
rect 1268 1137 1292 1143
rect 1316 1137 1420 1143
rect 1444 1137 1500 1143
rect 1524 1137 1676 1143
rect 1716 1137 2131 1143
rect 180 1117 220 1123
rect 740 1117 780 1123
rect 948 1117 956 1123
rect 980 1117 1084 1123
rect 1092 1117 1132 1123
rect 1252 1117 1308 1123
rect 1332 1117 1452 1123
rect 1540 1117 1644 1123
rect 1661 1117 1708 1123
rect 13 1104 19 1116
rect 212 1097 268 1103
rect 468 1097 524 1103
rect 532 1097 572 1103
rect 580 1097 588 1103
rect 612 1097 908 1103
rect 916 1097 1148 1103
rect 1156 1097 1196 1103
rect 1204 1097 1260 1103
rect 1268 1097 1388 1103
rect 1485 1103 1491 1116
rect 1661 1103 1667 1117
rect 1764 1117 1836 1123
rect 2125 1123 2131 1137
rect 2148 1137 2460 1143
rect 2596 1137 2620 1143
rect 2628 1137 2828 1143
rect 3028 1137 3052 1143
rect 3092 1137 3292 1143
rect 3316 1137 3372 1143
rect 3380 1137 3724 1143
rect 3732 1137 3788 1143
rect 3796 1137 4044 1143
rect 4052 1137 4076 1143
rect 4084 1137 4524 1143
rect 4564 1137 4796 1143
rect 4884 1137 4908 1143
rect 4948 1137 5004 1143
rect 5108 1137 5292 1143
rect 5357 1137 5484 1143
rect 1892 1117 1939 1123
rect 2125 1117 2172 1123
rect 1412 1097 1491 1103
rect 1517 1097 1667 1103
rect 84 1077 380 1083
rect 388 1077 428 1083
rect 468 1077 524 1083
rect 580 1077 915 1083
rect 52 1057 76 1063
rect 276 1057 300 1063
rect 500 1057 556 1063
rect 564 1057 620 1063
rect 628 1057 636 1063
rect 660 1057 668 1063
rect 724 1057 780 1063
rect 852 1057 876 1063
rect 909 1063 915 1077
rect 1108 1077 1164 1083
rect 1517 1083 1523 1097
rect 1684 1097 1740 1103
rect 1796 1097 1916 1103
rect 1933 1103 1939 1117
rect 2228 1117 2364 1123
rect 2372 1117 2412 1123
rect 2452 1117 2508 1123
rect 2532 1117 2540 1123
rect 2564 1117 2604 1123
rect 2756 1117 2940 1123
rect 2948 1117 3180 1123
rect 3268 1117 3516 1123
rect 3540 1117 3916 1123
rect 4180 1117 4332 1123
rect 4340 1117 4428 1123
rect 4468 1117 4524 1123
rect 4564 1117 4595 1123
rect 1933 1097 1948 1103
rect 2020 1097 2060 1103
rect 2132 1097 2604 1103
rect 2676 1097 3340 1103
rect 3380 1097 3532 1103
rect 3572 1097 3580 1103
rect 3764 1097 3852 1103
rect 3908 1097 4172 1103
rect 4308 1097 4364 1103
rect 4388 1097 4556 1103
rect 4589 1103 4595 1117
rect 4612 1117 4620 1123
rect 4660 1117 4748 1123
rect 4852 1117 5116 1123
rect 5140 1117 5180 1123
rect 5188 1117 5276 1123
rect 5357 1123 5363 1137
rect 5604 1137 5740 1143
rect 5780 1137 5836 1143
rect 5892 1137 5916 1143
rect 5972 1137 6012 1143
rect 6052 1137 6124 1143
rect 5284 1117 5363 1123
rect 5380 1117 5836 1123
rect 5853 1117 5868 1123
rect 4589 1097 4611 1103
rect 1492 1077 1523 1083
rect 1540 1077 1612 1083
rect 1652 1077 1708 1083
rect 1716 1077 1804 1083
rect 1860 1077 1868 1083
rect 1940 1077 2076 1083
rect 2164 1077 2188 1083
rect 2276 1077 2307 1083
rect 909 1057 1116 1063
rect 1156 1057 1564 1063
rect 1581 1057 1772 1063
rect 180 1037 316 1043
rect 356 1037 940 1043
rect 948 1037 1116 1043
rect 1124 1037 1260 1043
rect 1268 1037 1292 1043
rect 1581 1043 1587 1057
rect 1828 1057 1964 1063
rect 2020 1057 2060 1063
rect 2084 1057 2188 1063
rect 2212 1057 2220 1063
rect 2228 1057 2252 1063
rect 2260 1057 2268 1063
rect 2301 1063 2307 1077
rect 2324 1077 2444 1083
rect 2468 1077 2492 1083
rect 2548 1077 2732 1083
rect 2756 1077 2924 1083
rect 3108 1077 3244 1083
rect 3300 1077 3420 1083
rect 3524 1077 3532 1083
rect 3828 1077 4364 1083
rect 4436 1077 4588 1083
rect 4605 1083 4611 1097
rect 4628 1097 4732 1103
rect 4820 1097 4972 1103
rect 4996 1097 5372 1103
rect 5540 1097 5548 1103
rect 5588 1097 5628 1103
rect 5668 1097 5692 1103
rect 5716 1097 5788 1103
rect 5853 1103 5859 1117
rect 5892 1117 6108 1123
rect 6212 1117 6252 1123
rect 5805 1097 5859 1103
rect 5805 1084 5811 1097
rect 5876 1097 6220 1103
rect 4605 1077 4780 1083
rect 4884 1077 4972 1083
rect 5012 1077 5052 1083
rect 5076 1077 5100 1083
rect 5124 1077 5148 1083
rect 5316 1077 5324 1083
rect 5380 1077 5420 1083
rect 5524 1077 5532 1083
rect 5556 1077 5708 1083
rect 5732 1077 5772 1083
rect 5828 1077 5932 1083
rect 5972 1077 5980 1083
rect 6004 1077 6076 1083
rect 6100 1077 6124 1083
rect 6180 1077 6284 1083
rect 2301 1057 2428 1063
rect 2484 1057 2540 1063
rect 2644 1057 2892 1063
rect 2964 1057 3244 1063
rect 3300 1057 3884 1063
rect 4212 1057 4332 1063
rect 4388 1057 4844 1063
rect 4884 1057 5420 1063
rect 5444 1057 5484 1063
rect 5636 1057 5756 1063
rect 5876 1057 5964 1063
rect 6004 1057 6028 1063
rect 6084 1057 6108 1063
rect 6116 1057 6188 1063
rect 1364 1037 1587 1043
rect 1652 1037 1676 1043
rect 1716 1037 1731 1043
rect 100 1017 572 1023
rect 612 1017 988 1023
rect 1028 1017 1123 1023
rect 340 997 428 1003
rect 628 997 716 1003
rect 820 997 828 1003
rect 852 997 860 1003
rect 884 997 892 1003
rect 932 997 956 1003
rect 980 997 988 1003
rect 1076 997 1100 1003
rect 1117 1003 1123 1017
rect 1140 1017 1340 1023
rect 1380 1017 1516 1023
rect 1572 1017 1596 1023
rect 1684 1017 1708 1023
rect 1725 1023 1731 1037
rect 1789 1043 1795 1056
rect 1748 1037 1795 1043
rect 1860 1037 1916 1043
rect 1972 1037 2332 1043
rect 2388 1037 2460 1043
rect 2484 1037 2604 1043
rect 2628 1037 2764 1043
rect 2804 1037 2892 1043
rect 2932 1037 3068 1043
rect 3076 1037 3484 1043
rect 3556 1037 3596 1043
rect 3604 1037 3628 1043
rect 3668 1037 3916 1043
rect 4004 1037 4188 1043
rect 4212 1037 4332 1043
rect 4372 1037 4460 1043
rect 4484 1037 4652 1043
rect 4804 1037 4844 1043
rect 4852 1037 4988 1043
rect 4996 1037 5052 1043
rect 5060 1037 5228 1043
rect 5252 1037 5308 1043
rect 5332 1037 5372 1043
rect 5412 1037 5484 1043
rect 5508 1037 5612 1043
rect 5636 1037 5772 1043
rect 5828 1037 6044 1043
rect 1725 1017 1820 1023
rect 1908 1017 1980 1023
rect 2004 1017 2060 1023
rect 2100 1017 2156 1023
rect 2196 1017 2316 1023
rect 2356 1017 2380 1023
rect 2404 1017 2972 1023
rect 3028 1017 3084 1023
rect 3412 1017 3468 1023
rect 3492 1017 3804 1023
rect 3901 1017 4268 1023
rect 3112 1014 3160 1016
rect 3112 1006 3113 1014
rect 3122 1006 3123 1014
rect 3158 1006 3160 1014
rect 3112 1004 3160 1006
rect 1117 997 1164 1003
rect 1204 997 1388 1003
rect 1428 997 1516 1003
rect 1556 997 1756 1003
rect 1780 997 1964 1003
rect 2004 997 2220 1003
rect 2228 997 2236 1003
rect 2260 997 2332 1003
rect 2340 997 2396 1003
rect 2420 997 2540 1003
rect 2676 997 3084 1003
rect 3252 997 3491 1003
rect 132 977 204 983
rect 276 977 444 983
rect 740 977 940 983
rect 1028 977 1084 983
rect 1252 977 1372 983
rect 1460 977 1644 983
rect 1908 977 2044 983
rect 2084 977 2092 983
rect 2132 977 2316 983
rect 2420 977 2764 983
rect 2868 977 3036 983
rect 3252 977 3340 983
rect 3396 977 3420 983
rect 3485 983 3491 997
rect 3508 997 3516 1003
rect 3524 997 3612 1003
rect 3901 1003 3907 1017
rect 4372 1017 4540 1023
rect 4564 1017 4700 1023
rect 4788 1017 4972 1023
rect 4980 1017 5036 1023
rect 5044 1017 5068 1023
rect 5092 1017 5388 1023
rect 5524 1017 5564 1023
rect 5620 1017 5724 1023
rect 5844 1017 5868 1023
rect 6052 1017 6268 1023
rect 3652 997 3907 1003
rect 3924 997 4204 1003
rect 4340 997 4780 1003
rect 4852 997 5036 1003
rect 5172 997 5276 1003
rect 5284 997 5420 1003
rect 5428 997 5436 1003
rect 5444 997 5516 1003
rect 5620 997 5676 1003
rect 5860 997 6188 1003
rect 3485 977 3692 983
rect 3988 977 4124 983
rect 4164 977 4268 983
rect 4276 977 4316 983
rect 4500 977 4604 983
rect 4612 977 4620 983
rect 4820 977 4892 983
rect 4932 977 4988 983
rect 5028 977 5468 983
rect 5476 977 5836 983
rect 5844 977 5980 983
rect 6004 977 6028 983
rect 6180 980 6252 983
rect 6180 977 6259 980
rect 3373 964 3379 976
rect 148 957 172 963
rect 276 957 300 963
rect 308 957 364 963
rect 436 957 556 963
rect 692 957 716 963
rect 868 957 988 963
rect 1012 957 1068 963
rect 1092 957 1148 963
rect 1236 957 1292 963
rect 1396 957 1452 963
rect 1460 957 1468 963
rect 1492 957 1580 963
rect 1636 957 1676 963
rect 1732 957 1772 963
rect 1780 957 1836 963
rect 1844 957 1868 963
rect 1924 957 1948 963
rect 1988 957 1996 963
rect 2068 957 2108 963
rect 2116 957 2124 963
rect 2164 957 2220 963
rect 2276 957 2284 963
rect 2356 957 2412 963
rect 2436 957 2540 963
rect 2564 957 2588 963
rect 2660 957 2812 963
rect 2868 957 2972 963
rect 3076 957 3100 963
rect 3140 957 3276 963
rect 3396 957 3484 963
rect 3508 957 3564 963
rect 3604 957 3692 963
rect 3716 957 4108 963
rect 4196 957 4268 963
rect 4356 957 4428 963
rect 4468 957 5100 963
rect 5108 957 5132 963
rect 5156 957 5212 963
rect 5236 957 5324 963
rect 5364 957 5388 963
rect 5428 957 5516 963
rect 5540 957 5580 963
rect 5636 957 5660 963
rect 5700 957 5708 963
rect 5716 957 5740 963
rect 5844 957 5996 963
rect 6052 957 6108 963
rect 6212 957 6236 963
rect 20 937 140 943
rect 148 937 188 943
rect 260 937 300 943
rect 308 937 396 943
rect 484 937 524 943
rect 637 937 700 943
rect 212 917 316 923
rect 324 917 476 923
rect 637 923 643 937
rect 756 937 812 943
rect 884 937 1020 943
rect 1044 937 1052 943
rect 1076 937 1244 943
rect 1284 937 1308 943
rect 1316 937 1340 943
rect 1469 937 2172 943
rect 509 917 643 923
rect 509 903 515 917
rect 660 917 684 923
rect 692 917 700 923
rect 1469 923 1475 937
rect 2180 937 2444 943
rect 2452 937 2732 943
rect 2772 937 2828 943
rect 2868 937 2908 943
rect 2996 937 3004 943
rect 3220 937 3331 943
rect 708 917 1475 923
rect 1540 917 1628 923
rect 1764 917 1772 923
rect 1812 917 1836 923
rect 1844 917 1996 923
rect 2068 917 2092 923
rect 2180 917 2204 923
rect 2628 917 2668 923
rect 2676 917 2796 923
rect 2932 917 2988 923
rect 2996 917 3068 923
rect 3325 923 3331 937
rect 3348 937 3660 943
rect 3748 937 3836 943
rect 3908 937 3980 943
rect 4020 937 4908 943
rect 5012 937 5196 943
rect 5300 937 5324 943
rect 5348 937 5420 943
rect 5444 940 5484 943
rect 5444 937 5491 940
rect 5508 937 5596 943
rect 5620 937 5708 943
rect 5716 937 5724 943
rect 5812 937 5900 943
rect 5924 937 5932 943
rect 5940 937 5996 943
rect 6132 937 6236 943
rect 3204 917 3315 923
rect 3325 917 3500 923
rect 484 897 515 903
rect 525 897 652 903
rect 525 883 531 897
rect 660 897 796 903
rect 820 897 828 903
rect 916 897 972 903
rect 996 897 1116 903
rect 1396 897 1548 903
rect 1652 897 1692 903
rect 1716 897 1756 903
rect 1828 897 1868 903
rect 1892 897 2252 903
rect 2324 897 2524 903
rect 2548 897 2572 903
rect 2596 897 2860 903
rect 2932 897 2988 903
rect 3076 897 3212 903
rect 3220 897 3228 903
rect 3309 903 3315 917
rect 3556 917 3564 923
rect 4148 917 4220 923
rect 4228 917 4460 923
rect 4516 917 4572 923
rect 4628 917 4636 923
rect 4644 917 4732 923
rect 4749 917 4876 923
rect 3309 897 3340 903
rect 3476 897 3500 903
rect 3524 897 3708 903
rect 3828 897 3884 903
rect 4116 897 4188 903
rect 4228 897 4332 903
rect 4356 897 4396 903
rect 4420 897 4476 903
rect 4596 897 4620 903
rect 4749 903 4755 917
rect 4900 917 5020 923
rect 5060 917 5084 923
rect 5108 917 5164 923
rect 5220 917 5276 923
rect 5316 917 5452 923
rect 5476 920 5491 923
rect 5476 917 5484 920
rect 5508 917 5532 923
rect 5572 917 5603 923
rect 4644 897 4755 903
rect 4788 897 4812 903
rect 4884 897 5004 903
rect 5076 897 5228 903
rect 5268 897 5292 903
rect 5300 897 5436 903
rect 5469 897 5548 903
rect 1261 884 1267 896
rect 5069 884 5075 896
rect 5469 884 5475 897
rect 5597 903 5603 917
rect 5652 917 5676 923
rect 5732 917 5804 923
rect 5908 917 6252 923
rect 6292 917 6307 923
rect 5597 897 5763 903
rect 196 877 531 883
rect 564 877 668 883
rect 692 877 940 883
rect 964 877 1164 883
rect 1172 877 1212 883
rect 1300 877 1388 883
rect 1508 877 1516 883
rect 1556 877 2252 883
rect 2324 877 2860 883
rect 3028 877 3084 883
rect 3108 877 3196 883
rect 3316 877 3404 883
rect 3444 877 3676 883
rect 3693 877 4156 883
rect 260 857 508 863
rect 516 857 636 863
rect 676 857 972 863
rect 980 857 1100 863
rect 1124 857 1180 863
rect 1204 857 1340 863
rect 1380 857 1932 863
rect 1956 857 2012 863
rect 2052 857 2092 863
rect 2132 857 2252 863
rect 2292 857 2380 863
rect 2388 857 2428 863
rect 2452 857 2556 863
rect 2852 857 2908 863
rect 2948 857 2972 863
rect 3060 857 3532 863
rect 3556 857 3644 863
rect 3693 863 3699 877
rect 4196 877 4236 883
rect 4244 877 4284 883
rect 4308 877 4348 883
rect 4436 877 4540 883
rect 4564 877 4668 883
rect 4772 877 4892 883
rect 4916 877 4956 883
rect 4980 877 5020 883
rect 5124 877 5244 883
rect 5332 877 5388 883
rect 5492 877 5548 883
rect 5556 877 5740 883
rect 5757 883 5763 897
rect 5796 897 5932 903
rect 6084 897 6108 903
rect 6164 897 6284 903
rect 5757 877 5836 883
rect 5892 877 5900 883
rect 6036 877 6060 883
rect 6068 877 6076 883
rect 6301 883 6307 917
rect 6260 877 6307 883
rect 3668 857 3699 863
rect 3860 857 4940 863
rect 4948 857 5356 863
rect 5396 857 5436 863
rect 5460 857 5516 863
rect 5572 857 5612 863
rect 5636 857 5660 863
rect 5684 860 5772 863
rect 5684 857 5779 860
rect 5892 857 5932 863
rect 6004 857 6252 863
rect 637 837 748 843
rect 324 817 348 823
rect 436 817 492 823
rect 637 823 643 837
rect 788 837 1324 843
rect 1332 837 2348 843
rect 2404 837 2412 843
rect 2484 837 2636 843
rect 2660 837 3100 843
rect 3124 837 3244 843
rect 3252 837 3308 843
rect 3348 837 3500 843
rect 3524 837 3564 843
rect 3588 837 4108 843
rect 4148 837 4588 843
rect 4596 837 5052 843
rect 5076 837 5628 843
rect 5636 837 5676 843
rect 5700 840 5779 843
rect 5700 837 5772 840
rect 5972 837 6236 843
rect 6244 837 6284 843
rect 516 817 643 823
rect 756 817 780 823
rect 820 817 1052 823
rect 1380 817 1548 823
rect 1748 817 2044 823
rect 2052 817 2124 823
rect 2148 817 2188 823
rect 2196 817 2284 823
rect 2292 817 2332 823
rect 2356 817 2940 823
rect 2948 817 3852 823
rect 3924 817 3996 823
rect 4036 817 4323 823
rect 1576 814 1624 816
rect 1576 806 1577 814
rect 1586 806 1587 814
rect 1622 806 1624 814
rect 1576 804 1624 806
rect 340 797 364 803
rect 372 797 764 803
rect 772 797 1036 803
rect 1044 797 1100 803
rect 1108 797 1196 803
rect 1204 797 1244 803
rect 1428 797 1468 803
rect 1476 797 1555 803
rect 468 777 716 783
rect 772 777 812 783
rect 948 777 1068 783
rect 1140 777 1388 783
rect 1549 783 1555 797
rect 1748 797 1916 803
rect 2068 797 2156 803
rect 2164 797 2284 803
rect 2308 797 2764 803
rect 2788 797 2812 803
rect 2852 797 3020 803
rect 3060 797 3068 803
rect 3092 797 3740 803
rect 3892 797 4300 803
rect 4317 803 4323 817
rect 4340 817 4364 823
rect 4372 817 4412 823
rect 4436 817 4508 823
rect 4580 817 4588 823
rect 4756 817 5068 823
rect 5092 817 5132 823
rect 5156 817 5308 823
rect 5332 817 5420 823
rect 5444 817 5644 823
rect 5812 817 5852 823
rect 5892 817 5980 823
rect 6052 817 6284 823
rect 4664 814 4712 816
rect 4664 806 4665 814
rect 4674 806 4675 814
rect 4710 806 4712 814
rect 4664 804 4712 806
rect 4317 797 4332 803
rect 4388 797 4396 803
rect 4404 797 4460 803
rect 4500 797 4524 803
rect 4756 797 4956 803
rect 4980 797 5724 803
rect 5732 797 6076 803
rect 1549 777 1900 783
rect 1908 777 2508 783
rect 2548 777 2716 783
rect 2996 777 3596 783
rect 3604 777 3660 783
rect 3876 777 4444 783
rect 4500 777 4668 783
rect 4676 777 4908 783
rect 4916 777 4940 783
rect 5076 777 5260 783
rect 5284 777 5331 783
rect 916 757 1084 763
rect 1108 757 1148 763
rect 1188 757 1388 763
rect 1444 757 1452 763
rect 1540 757 1596 763
rect 1652 757 1836 763
rect 1876 757 1948 763
rect 2036 757 2124 763
rect 2141 757 2172 763
rect 68 737 716 743
rect 724 737 1116 743
rect 1124 737 1276 743
rect 1332 737 1340 743
rect 1444 737 1468 743
rect 1492 737 1580 743
rect 1652 737 1692 743
rect 1741 737 1884 743
rect 452 717 524 723
rect 532 717 540 723
rect 596 717 620 723
rect 644 717 684 723
rect 692 717 780 723
rect 820 717 828 723
rect 980 717 1043 723
rect 452 697 492 703
rect 996 697 1020 703
rect 1037 684 1043 717
rect 1741 723 1747 737
rect 1940 737 1964 743
rect 2004 737 2060 743
rect 2141 743 2147 757
rect 2212 757 2236 763
rect 2260 757 2284 763
rect 2308 757 2476 763
rect 2500 757 2764 763
rect 2836 757 3340 763
rect 3428 757 3580 763
rect 3620 757 3820 763
rect 4116 757 4828 763
rect 4836 757 4940 763
rect 5012 757 5068 763
rect 5108 757 5132 763
rect 5172 757 5276 763
rect 5325 763 5331 777
rect 5364 777 5372 783
rect 5476 777 5596 783
rect 5620 777 5692 783
rect 5716 777 5916 783
rect 5972 777 6012 783
rect 6068 777 6124 783
rect 5325 757 5468 763
rect 5540 757 5740 763
rect 5812 757 5836 763
rect 5908 757 6092 763
rect 6100 757 6252 763
rect 2068 737 2147 743
rect 2196 737 2204 743
rect 2228 737 2275 743
rect 1060 717 1747 723
rect 1764 717 1852 723
rect 1876 717 2124 723
rect 2196 717 2252 723
rect 2269 723 2275 737
rect 2324 737 2444 743
rect 2468 737 2524 743
rect 2580 737 2604 743
rect 2612 737 2828 743
rect 3012 737 3020 743
rect 3476 737 3484 743
rect 3508 737 3699 743
rect 2269 717 2572 723
rect 2596 717 2604 723
rect 2644 717 2828 723
rect 2916 717 3244 723
rect 3268 717 3276 723
rect 3316 717 3372 723
rect 3412 717 3516 723
rect 3620 717 3676 723
rect 3693 723 3699 737
rect 4212 737 4732 743
rect 4740 737 5100 743
rect 5108 737 5484 743
rect 5492 737 6060 743
rect 6093 737 6156 743
rect 3693 717 3916 723
rect 4068 717 4092 723
rect 4148 717 4204 723
rect 4308 717 4332 723
rect 4356 717 4428 723
rect 4436 717 4460 723
rect 4500 717 4604 723
rect 4628 717 4748 723
rect 4772 717 4828 723
rect 4980 717 5004 723
rect 5028 717 5148 723
rect 5844 717 5932 723
rect 6093 723 6099 737
rect 6244 737 6284 743
rect 6061 717 6099 723
rect 1060 700 1132 703
rect 2157 704 2163 716
rect 1140 700 1260 703
rect 1060 697 1260 700
rect 1300 697 1756 703
rect 1876 697 2019 703
rect 52 677 124 683
rect 228 677 332 683
rect 340 677 348 683
rect 580 677 620 683
rect 628 677 892 683
rect 900 677 908 683
rect 964 677 1004 683
rect 1092 677 1116 683
rect 1133 680 1164 683
rect 1140 677 1164 680
rect 1268 677 1324 683
rect 1332 677 1372 683
rect 1476 677 1548 683
rect 2013 683 2019 697
rect 2036 697 2092 703
rect 2100 697 2156 703
rect 2180 697 2444 703
rect 2468 697 2684 703
rect 2692 697 2755 703
rect 2013 677 2028 683
rect 2052 677 2172 683
rect 2196 677 2236 683
rect 2244 677 2396 683
rect 2420 677 2444 683
rect 2541 677 2652 683
rect 20 657 60 663
rect 68 657 140 663
rect 148 657 204 663
rect 612 657 972 663
rect 1076 657 1132 663
rect 1172 657 1228 663
rect 1268 657 1740 663
rect 1780 657 1948 663
rect 1956 657 2060 663
rect 2116 657 2131 663
rect 356 637 428 643
rect 436 637 476 643
rect 484 637 524 643
rect 564 637 748 643
rect 1108 640 1164 643
rect 1108 637 1171 640
rect 1268 637 1484 643
rect 1540 637 1660 643
rect 1668 637 1724 643
rect 1732 637 1740 643
rect 1764 637 2108 643
rect 2125 643 2131 657
rect 2164 657 2259 663
rect 2125 637 2172 643
rect 2196 637 2220 643
rect 2253 643 2259 657
rect 2276 657 2332 663
rect 2541 663 2547 677
rect 2676 677 2700 683
rect 2749 683 2755 697
rect 2932 697 2972 703
rect 2989 697 3196 703
rect 2749 677 2780 683
rect 2989 683 2995 697
rect 3220 697 3292 703
rect 3444 697 3628 703
rect 3636 697 3644 703
rect 3828 697 3900 703
rect 3988 697 4028 703
rect 4052 697 4220 703
rect 4308 697 4883 703
rect 2836 677 2995 683
rect 3076 677 3132 683
rect 3316 677 3436 683
rect 3444 677 3468 683
rect 3725 683 3731 696
rect 3524 677 3788 683
rect 3812 677 4012 683
rect 4164 677 4204 683
rect 4276 677 4364 683
rect 4388 677 4556 683
rect 4596 677 4604 683
rect 4612 677 4748 683
rect 4772 677 4812 683
rect 4877 683 4883 697
rect 5204 697 5244 703
rect 5268 697 5356 703
rect 5492 697 5500 703
rect 5524 697 5667 703
rect 4877 677 5308 683
rect 5661 683 5667 697
rect 5700 697 5788 703
rect 5796 697 5820 703
rect 5828 697 5852 703
rect 6061 703 6067 717
rect 6116 717 6156 723
rect 6253 704 6259 716
rect 6020 697 6067 703
rect 6084 697 6195 703
rect 5348 677 5651 683
rect 5661 677 5900 683
rect 2340 657 2547 663
rect 2564 657 2668 663
rect 2772 657 2812 663
rect 2820 657 2972 663
rect 3108 657 3148 663
rect 3252 657 3612 663
rect 3748 657 3756 663
rect 3764 657 3852 663
rect 3860 657 4108 663
rect 4125 657 4412 663
rect 2253 637 2524 643
rect 2548 637 2572 643
rect 2596 637 2780 643
rect 2804 637 2956 643
rect 2980 637 3052 643
rect 3060 637 3228 643
rect 3236 637 3324 643
rect 3332 637 3548 643
rect 3588 637 3836 643
rect 3844 637 4028 643
rect 4125 643 4131 657
rect 4580 657 4723 663
rect 4100 637 4131 643
rect 4164 637 4220 643
rect 4253 637 4483 643
rect 116 617 444 623
rect 468 617 508 623
rect 564 617 812 623
rect 820 617 844 623
rect 852 617 940 623
rect 964 617 988 623
rect 1044 617 1132 623
rect 1165 620 1276 623
rect 1172 617 1276 620
rect 1668 617 1836 623
rect 1860 617 1868 623
rect 1876 617 1932 623
rect 1972 617 1996 623
rect 2052 617 2060 623
rect 2132 617 2556 623
rect 2580 617 2588 623
rect 2596 617 2668 623
rect 2708 617 2860 623
rect 2868 617 2892 623
rect 2932 617 3020 623
rect 3236 617 3244 623
rect 3268 617 3436 623
rect 3460 617 3484 623
rect 3501 617 3996 623
rect 3112 614 3160 616
rect 3112 606 3113 614
rect 3122 606 3123 614
rect 3158 606 3160 614
rect 3112 604 3160 606
rect 388 597 1116 603
rect 1460 597 1875 603
rect 420 577 716 583
rect 804 577 979 583
rect 180 557 364 563
rect 452 557 588 563
rect 596 557 636 563
rect 660 557 732 563
rect 756 557 812 563
rect 836 557 908 563
rect 932 557 956 563
rect 973 563 979 577
rect 996 577 1052 583
rect 1060 577 1196 583
rect 1204 577 1324 583
rect 1332 577 1388 583
rect 1444 577 1516 583
rect 1556 577 1660 583
rect 1732 577 1740 583
rect 1869 583 1875 597
rect 1892 597 1964 603
rect 1972 597 1980 603
rect 1988 597 2108 603
rect 2116 597 2124 603
rect 2132 597 2236 603
rect 2260 597 2380 603
rect 2420 597 2588 603
rect 2628 597 2876 603
rect 2884 597 3091 603
rect 1869 577 2124 583
rect 2132 577 2364 583
rect 2452 577 2604 583
rect 2804 577 2844 583
rect 3085 583 3091 597
rect 3188 597 3372 603
rect 3501 603 3507 617
rect 4253 623 4259 637
rect 4020 617 4259 623
rect 4276 617 4332 623
rect 4340 617 4428 623
rect 4477 623 4483 637
rect 4532 637 4572 643
rect 4596 637 4652 643
rect 4717 643 4723 657
rect 4820 657 4972 663
rect 5156 657 5228 663
rect 5252 657 5292 663
rect 5332 657 5340 663
rect 5428 657 5452 663
rect 5460 657 5564 663
rect 5645 663 5651 677
rect 6004 677 6156 683
rect 6189 683 6195 697
rect 6189 677 6204 683
rect 6228 677 6252 683
rect 5645 657 5788 663
rect 5892 657 5948 663
rect 5972 657 5996 663
rect 6004 657 6060 663
rect 6100 657 6124 663
rect 4717 637 4764 643
rect 4788 637 4876 643
rect 4884 637 4924 643
rect 4964 637 5052 643
rect 5364 637 5596 643
rect 5604 637 5644 643
rect 5652 637 5676 643
rect 5764 637 5916 643
rect 6132 637 6252 643
rect 4477 617 4620 623
rect 4884 617 4940 623
rect 5012 617 5228 623
rect 5268 617 5356 623
rect 5380 617 5388 623
rect 5428 617 5468 623
rect 5556 617 5628 623
rect 6116 617 6220 623
rect 3396 597 3507 603
rect 3524 597 3644 603
rect 3748 597 3772 603
rect 3796 597 3884 603
rect 4004 597 4140 603
rect 4420 597 4972 603
rect 4980 597 4988 603
rect 5044 597 5068 603
rect 5124 597 5212 603
rect 5236 597 5260 603
rect 5348 597 5516 603
rect 5572 597 5676 603
rect 5748 597 5827 603
rect 3085 577 3116 583
rect 3172 577 3228 583
rect 3284 577 3628 583
rect 3796 577 3836 583
rect 3876 577 3948 583
rect 3988 577 4156 583
rect 4308 577 4419 583
rect 3661 564 3667 576
rect 973 557 1628 563
rect 1636 557 1996 563
rect 2013 557 2076 563
rect 500 537 556 543
rect 564 537 572 543
rect 628 537 652 543
rect 676 537 860 543
rect 925 537 1100 543
rect 260 517 492 523
rect 692 517 700 523
rect 925 523 931 537
rect 1140 537 1148 543
rect 1332 537 1372 543
rect 1412 537 1468 543
rect 1492 537 1644 543
rect 1684 537 1692 543
rect 1700 537 1724 543
rect 1748 537 1772 543
rect 1821 537 1868 543
rect 756 517 931 523
rect 1044 517 1436 523
rect 1460 517 1500 523
rect 1508 517 1532 523
rect 1604 517 1763 523
rect 941 504 947 516
rect 148 497 556 503
rect 596 497 780 503
rect 788 497 812 503
rect 964 497 1116 503
rect 1156 497 1324 503
rect 1412 497 1484 503
rect 1684 497 1708 503
rect 1757 503 1763 517
rect 1821 503 1827 537
rect 2013 543 2019 557
rect 2100 557 2156 563
rect 2196 557 2364 563
rect 2388 557 2620 563
rect 2772 557 2860 563
rect 3076 557 3132 563
rect 3220 557 3228 563
rect 3300 557 3308 563
rect 3380 557 3564 563
rect 3588 557 3628 563
rect 3684 557 3740 563
rect 3764 557 3788 563
rect 3828 557 3916 563
rect 3924 557 3980 563
rect 4020 557 4108 563
rect 4180 557 4204 563
rect 4292 557 4316 563
rect 4413 563 4419 577
rect 4436 577 4460 583
rect 4500 577 4524 583
rect 4541 577 4652 583
rect 4541 563 4547 577
rect 4660 577 4796 583
rect 4820 577 4908 583
rect 4932 577 4940 583
rect 5012 577 5164 583
rect 5204 577 5420 583
rect 5780 577 5804 583
rect 5821 583 5827 597
rect 5844 597 5868 603
rect 5892 597 5932 603
rect 6004 597 6284 603
rect 5821 577 5948 583
rect 6004 577 6140 583
rect 4413 557 4547 563
rect 4756 560 4876 563
rect 4749 557 4876 560
rect 5108 557 5260 563
rect 5300 557 5372 563
rect 5405 557 5516 563
rect 1908 537 2019 543
rect 2036 537 2172 543
rect 2212 537 2252 543
rect 2260 537 2316 543
rect 2388 537 2476 543
rect 2484 537 2524 543
rect 2621 537 2636 543
rect 1837 517 1932 523
rect 1837 504 1843 517
rect 1972 517 2188 523
rect 2228 517 2284 523
rect 2308 517 2348 523
rect 2372 517 2412 523
rect 2436 517 2572 523
rect 2621 523 2627 537
rect 2676 537 2748 543
rect 2756 537 2780 543
rect 2964 537 2988 543
rect 3108 537 3324 543
rect 3348 537 3420 543
rect 3540 537 3596 543
rect 3748 537 3804 543
rect 3828 537 4012 543
rect 4036 537 4060 543
rect 4132 537 4140 543
rect 4276 537 4604 543
rect 4628 540 4755 543
rect 4628 537 4748 540
rect 2596 517 2627 523
rect 2740 517 2748 523
rect 2829 523 2835 536
rect 4820 537 5228 543
rect 5405 543 5411 557
rect 5556 557 5804 563
rect 5812 557 5916 563
rect 5869 544 5875 557
rect 5940 557 6060 563
rect 6084 557 6140 563
rect 6164 557 6204 563
rect 6260 557 6284 563
rect 5268 537 5411 543
rect 5428 537 5484 543
rect 5588 537 5708 543
rect 5844 537 5852 543
rect 5972 537 6252 543
rect 2829 517 2860 523
rect 2916 517 2972 523
rect 2996 517 3020 523
rect 3044 517 3084 523
rect 3124 517 3324 523
rect 3348 517 3356 523
rect 3380 517 3436 523
rect 3524 517 3747 523
rect 2637 504 2643 516
rect 1757 497 1827 503
rect 1860 497 1916 503
rect 1956 497 2140 503
rect 2164 497 2220 503
rect 2228 497 2492 503
rect 2500 497 2572 503
rect 2660 497 2764 503
rect 2820 497 2828 503
rect 2852 497 2924 503
rect 2932 497 3020 503
rect 3060 497 3068 503
rect 3508 497 3692 503
rect 3716 497 3724 503
rect 3741 503 3747 517
rect 3780 517 3788 523
rect 3924 517 4300 523
rect 4356 517 4460 523
rect 4500 517 4540 523
rect 4548 517 4796 523
rect 4820 517 4908 523
rect 4932 517 5004 523
rect 5076 517 5084 523
rect 5124 517 5132 523
rect 5188 517 5244 523
rect 5252 517 5420 523
rect 5549 523 5555 536
rect 5460 517 5612 523
rect 5636 517 5916 523
rect 6100 517 6284 523
rect 3741 497 3868 503
rect 3940 497 3964 503
rect 3981 497 4236 503
rect 20 477 604 483
rect 612 477 620 483
rect 644 477 748 483
rect 772 477 844 483
rect 1204 477 2540 483
rect 2548 477 2796 483
rect 2900 477 3452 483
rect 3981 483 3987 497
rect 4260 497 4268 503
rect 4340 497 4492 503
rect 4564 497 4700 503
rect 4756 497 4860 503
rect 4884 497 4988 503
rect 5005 503 5011 516
rect 5005 497 5356 503
rect 5364 497 5388 503
rect 5444 497 5468 503
rect 5476 497 5500 503
rect 5556 497 5868 503
rect 5972 497 5996 503
rect 6020 497 6268 503
rect 3476 477 3987 483
rect 4020 477 4140 483
rect 4148 477 4268 483
rect 4292 477 4428 483
rect 4452 477 4908 483
rect 4916 477 5212 483
rect 5236 477 5340 483
rect 5428 477 5500 483
rect 5524 477 5596 483
rect 5620 477 5740 483
rect 5796 477 5996 483
rect 6148 477 6204 483
rect 1620 457 1932 463
rect 1940 457 1980 463
rect 2020 457 2044 463
rect 2068 457 2204 463
rect 2228 457 2316 463
rect 2340 457 3196 463
rect 3236 457 3260 463
rect 3284 457 3964 463
rect 4180 457 4588 463
rect 4708 457 4940 463
rect 4980 457 5020 463
rect 5044 457 5132 463
rect 5236 457 5276 463
rect 5332 457 5356 463
rect 5428 457 5564 463
rect 5588 457 5644 463
rect 5972 457 6076 463
rect 1556 437 1580 443
rect 1860 437 1884 443
rect 1940 437 2124 443
rect 2148 437 2460 443
rect 2484 437 2556 443
rect 2612 437 3756 443
rect 3773 437 3788 443
rect 740 417 844 423
rect 852 417 1084 423
rect 1092 417 1164 423
rect 1188 417 1516 423
rect 1725 417 1795 423
rect 1576 414 1624 416
rect 1576 406 1577 414
rect 1586 406 1587 414
rect 1622 406 1624 414
rect 1576 404 1624 406
rect 596 397 828 403
rect 884 397 1228 403
rect 1332 397 1404 403
rect 1428 397 1484 403
rect 1725 403 1731 417
rect 1652 397 1731 403
rect 1748 397 1772 403
rect 1789 403 1795 417
rect 1812 417 2140 423
rect 2164 417 2236 423
rect 2260 417 2316 423
rect 2324 417 2748 423
rect 2772 417 2924 423
rect 2932 417 3708 423
rect 3773 423 3779 437
rect 3860 437 3932 443
rect 3956 437 4044 443
rect 4068 437 4364 443
rect 4516 437 4636 443
rect 4692 437 6092 443
rect 3732 417 3779 423
rect 3908 417 4316 423
rect 4404 417 4579 423
rect 1789 397 1868 403
rect 1892 397 2396 403
rect 2420 397 2892 403
rect 2916 397 2956 403
rect 2980 397 2988 403
rect 3028 397 3148 403
rect 3252 397 3820 403
rect 3828 397 3900 403
rect 4020 397 4220 403
rect 4244 397 4476 403
rect 4573 403 4579 417
rect 4900 417 4972 423
rect 5044 417 5340 423
rect 5364 417 5452 423
rect 5508 417 5548 423
rect 5604 417 5772 423
rect 5805 417 6220 423
rect 4664 414 4712 416
rect 4664 406 4665 414
rect 4674 406 4675 414
rect 4710 406 4712 414
rect 4664 404 4712 406
rect 4573 397 4604 403
rect 4740 397 4796 403
rect 4868 397 4876 403
rect 4964 397 5036 403
rect 5156 397 5484 403
rect 5524 397 5692 403
rect 5805 403 5811 417
rect 5716 397 5811 403
rect 5940 397 5980 403
rect 6036 397 6108 403
rect 148 377 380 383
rect 1092 377 1132 383
rect 1140 377 1148 383
rect 1236 377 3324 383
rect 3348 377 3484 383
rect 3604 377 3612 383
rect 3700 377 3724 383
rect 3741 377 3916 383
rect 580 357 1539 363
rect 1060 337 1068 343
rect 1076 337 1260 343
rect 1268 337 1452 343
rect 1460 337 1516 343
rect 1533 343 1539 357
rect 1588 357 1932 363
rect 1972 357 2412 363
rect 2468 357 2716 363
rect 2804 357 3180 363
rect 3741 363 3747 377
rect 3940 377 4060 383
rect 4077 377 4204 383
rect 3188 357 3747 363
rect 3764 357 3788 363
rect 3812 357 3852 363
rect 3892 357 4028 363
rect 4077 363 4083 377
rect 4244 377 4604 383
rect 4756 377 4812 383
rect 4836 377 5091 383
rect 5085 364 5091 377
rect 5108 377 5164 383
rect 5204 377 5228 383
rect 5236 377 5676 383
rect 5732 377 5964 383
rect 5972 377 6172 383
rect 4052 357 4083 363
rect 4100 357 4156 363
rect 4180 357 4268 363
rect 4340 357 4460 363
rect 4468 357 4556 363
rect 4564 357 4620 363
rect 4628 357 4844 363
rect 4852 357 5068 363
rect 5092 357 5260 363
rect 5380 357 5468 363
rect 5492 357 5532 363
rect 5588 357 5772 363
rect 5796 357 5852 363
rect 5940 357 6012 363
rect 6045 357 6092 363
rect 1533 337 1596 343
rect 1652 337 2188 343
rect 2244 337 2332 343
rect 2349 337 2508 343
rect 884 317 1084 323
rect 1108 317 1180 323
rect 1204 317 1324 323
rect 1412 317 1500 323
rect 1508 317 1564 323
rect 1572 317 1628 323
rect 1668 317 1715 323
rect 84 297 108 303
rect 324 297 460 303
rect 468 297 492 303
rect 692 297 812 303
rect 1156 297 1276 303
rect 1300 300 1532 303
rect 1293 297 1532 300
rect 1556 297 1692 303
rect 1709 303 1715 317
rect 1732 317 1884 323
rect 1908 317 2156 323
rect 2164 317 2236 323
rect 2349 323 2355 337
rect 2580 337 2620 343
rect 2644 337 2668 343
rect 2740 337 2819 343
rect 2317 317 2355 323
rect 1709 297 1868 303
rect 2004 297 2028 303
rect 2100 297 2156 303
rect 2317 303 2323 317
rect 2372 317 2492 323
rect 2548 317 2604 323
rect 2644 317 2668 323
rect 2765 304 2771 316
rect 2196 297 2323 303
rect 2340 297 2348 303
rect 2372 297 2412 303
rect 2516 297 2620 303
rect 2637 297 2748 303
rect 1901 284 1907 296
rect 228 277 236 283
rect 724 277 924 283
rect 1220 277 1260 283
rect 1293 280 1308 283
rect 1300 277 1308 280
rect 1316 277 1324 283
rect 1348 277 1356 283
rect 1412 277 1420 283
rect 1492 277 1500 283
rect 1524 277 1612 283
rect 1748 277 1772 283
rect 1796 277 1884 283
rect 1940 277 2547 283
rect 196 257 364 263
rect 372 257 540 263
rect 548 257 892 263
rect 996 257 1228 263
rect 1316 257 1388 263
rect 1444 257 1724 263
rect 1732 257 1996 263
rect 2004 257 2060 263
rect 2084 257 2524 263
rect 2541 263 2547 277
rect 2637 283 2643 297
rect 2813 303 2819 337
rect 2884 337 2940 343
rect 2980 337 3196 343
rect 3220 337 3228 343
rect 3252 337 3292 343
rect 3332 337 3420 343
rect 3444 337 3532 343
rect 3556 337 3564 343
rect 3588 337 3612 343
rect 3668 337 3676 343
rect 3700 337 4188 343
rect 4196 337 4428 343
rect 4436 337 4492 343
rect 4500 337 4540 343
rect 4612 337 4732 343
rect 4788 337 5052 343
rect 5060 337 5276 343
rect 5284 337 5404 343
rect 5421 337 5676 343
rect 2957 324 2963 336
rect 2836 317 2860 323
rect 2996 317 3132 323
rect 3204 317 3516 323
rect 3540 317 3628 323
rect 3652 317 3708 323
rect 3732 317 3852 323
rect 3876 317 4236 323
rect 4276 317 4499 323
rect 2925 304 2931 316
rect 2813 297 2908 303
rect 2996 297 3715 303
rect 2612 277 2643 283
rect 2724 277 2908 283
rect 2932 277 2972 283
rect 2980 277 3068 283
rect 3092 277 3228 283
rect 3284 277 3324 283
rect 3348 277 3372 283
rect 3412 277 3436 283
rect 3492 277 3596 283
rect 3636 277 3692 283
rect 3709 283 3715 297
rect 3732 297 4092 303
rect 4116 297 4195 303
rect 3709 277 3916 283
rect 3940 277 4060 283
rect 4116 277 4140 283
rect 4189 283 4195 297
rect 4212 297 4476 303
rect 4493 303 4499 317
rect 4516 317 4524 323
rect 4564 317 4588 323
rect 4628 317 5004 323
rect 5012 317 5068 323
rect 5124 317 5180 323
rect 5188 317 5212 323
rect 5341 317 5356 323
rect 4493 297 4780 303
rect 4797 297 4812 303
rect 4189 277 4252 283
rect 4308 277 4364 283
rect 4404 277 4556 283
rect 4596 277 4707 283
rect 2541 257 2988 263
rect 3060 257 3484 263
rect 3524 257 3532 263
rect 3572 257 3660 263
rect 3668 257 3788 263
rect 3812 257 3836 263
rect 3860 257 3884 263
rect 3908 257 4076 263
rect 4084 257 4428 263
rect 4436 257 4460 263
rect 4500 257 4588 263
rect 4701 263 4707 277
rect 4797 283 4803 297
rect 4836 297 4876 303
rect 4884 297 4956 303
rect 5012 297 5020 303
rect 5108 297 5132 303
rect 5341 303 5347 317
rect 5421 323 5427 337
rect 5732 337 5788 343
rect 5940 337 6012 343
rect 5380 317 5427 323
rect 5437 317 5532 323
rect 5149 297 5347 303
rect 4772 277 4803 283
rect 5149 283 5155 297
rect 5437 303 5443 317
rect 5540 317 5580 323
rect 5668 317 5708 323
rect 5780 317 5852 323
rect 6045 323 6051 357
rect 6164 357 6188 363
rect 6061 324 6067 336
rect 5892 317 6051 323
rect 6077 317 6140 323
rect 5364 297 5443 303
rect 5476 297 5843 303
rect 4868 277 5155 283
rect 5172 277 5436 283
rect 5652 277 5676 283
rect 5780 277 5804 283
rect 5837 283 5843 297
rect 5860 297 5868 303
rect 5956 297 5964 303
rect 6077 303 6083 317
rect 6068 297 6083 303
rect 5837 277 5955 283
rect 4701 257 4844 263
rect 4852 257 4940 263
rect 4964 257 5020 263
rect 5044 257 5116 263
rect 5172 257 5420 263
rect 5460 257 5500 263
rect 5524 257 5932 263
rect 5949 263 5955 277
rect 5972 277 5996 283
rect 6100 277 6124 283
rect 5949 257 6028 263
rect 6052 257 6108 263
rect 6116 257 6252 263
rect 980 237 1084 243
rect 1124 237 1324 243
rect 1364 237 1532 243
rect 1556 237 1580 243
rect 1604 237 1964 243
rect 2020 237 2124 243
rect 2164 237 2204 243
rect 2260 237 2828 243
rect 2900 237 2940 243
rect 2964 237 3340 243
rect 3348 237 3948 243
rect 3956 237 4140 243
rect 4244 237 4332 243
rect 4340 237 4451 243
rect 660 217 876 223
rect 980 217 1660 223
rect 1684 217 1692 223
rect 1716 217 1884 223
rect 1908 217 1916 223
rect 1940 217 1964 223
rect 1988 217 2339 223
rect 1060 197 1196 203
rect 1252 197 1276 203
rect 1300 197 1340 203
rect 1364 197 1500 203
rect 1524 197 1740 203
rect 1780 197 1820 203
rect 1844 197 2044 203
rect 2052 197 2156 203
rect 2180 197 2316 203
rect 2333 203 2339 217
rect 2388 217 2396 223
rect 2420 217 2556 223
rect 2580 217 2668 223
rect 2692 217 2812 223
rect 2836 217 3052 223
rect 3204 217 3299 223
rect 3112 214 3160 216
rect 3112 206 3113 214
rect 3122 206 3123 214
rect 3158 206 3160 214
rect 3112 204 3160 206
rect 2333 197 2764 203
rect 2788 197 2796 203
rect 2820 197 2892 203
rect 2916 197 3004 203
rect 3012 197 3084 203
rect 3236 197 3244 203
rect 3293 203 3299 217
rect 3332 217 3420 223
rect 3460 217 3564 223
rect 3604 217 3724 223
rect 3748 217 3964 223
rect 3988 217 4028 223
rect 4036 217 4380 223
rect 4445 223 4451 237
rect 4468 237 4492 243
rect 4500 237 4604 243
rect 4644 237 4748 243
rect 4820 237 4988 243
rect 4996 237 5196 243
rect 5204 237 5228 243
rect 5236 237 5244 243
rect 5284 237 6156 243
rect 6164 237 6236 243
rect 4445 217 4588 223
rect 4692 217 4764 223
rect 4788 217 4876 223
rect 4980 217 5036 223
rect 5044 217 5340 223
rect 5348 217 6044 223
rect 6084 217 6156 223
rect 3293 197 3708 203
rect 3780 197 4524 203
rect 4532 197 4604 203
rect 4612 197 4668 203
rect 4676 197 4812 203
rect 4884 197 5203 203
rect 333 184 339 196
rect 772 177 780 183
rect 932 177 1068 183
rect 1076 177 1164 183
rect 1188 177 1708 183
rect 1732 177 1964 183
rect 1988 177 2028 183
rect 2068 177 2083 183
rect 852 157 860 163
rect 1076 157 1084 163
rect 1101 157 1260 163
rect 788 137 924 143
rect 1101 143 1107 157
rect 1277 157 1292 163
rect 1012 137 1107 143
rect 1277 143 1283 157
rect 1309 157 1356 163
rect 1172 137 1283 143
rect 1309 143 1315 157
rect 1396 157 1484 163
rect 1492 157 2060 163
rect 2077 163 2083 177
rect 2100 177 2316 183
rect 2356 177 2412 183
rect 2436 177 2540 183
rect 2548 177 3244 183
rect 3268 177 3276 183
rect 3316 177 3660 183
rect 3677 177 4108 183
rect 2077 157 2092 163
rect 2116 157 2195 163
rect 1300 137 1315 143
rect 1332 137 1372 143
rect 1380 137 2060 143
rect 2068 137 2140 143
rect 2189 143 2195 157
rect 2212 157 2252 163
rect 2308 157 2332 163
rect 2340 157 2428 163
rect 2468 157 2828 163
rect 2836 157 2956 163
rect 2980 157 3308 163
rect 3348 157 3468 163
rect 3492 157 3500 163
rect 3677 163 3683 177
rect 4148 177 4220 183
rect 4237 177 4380 183
rect 3540 157 3683 163
rect 3716 157 3804 163
rect 3924 157 4156 163
rect 4237 163 4243 177
rect 4397 177 4556 183
rect 4196 157 4243 163
rect 4276 157 4332 163
rect 4397 163 4403 177
rect 4628 177 5020 183
rect 5028 177 5036 183
rect 5092 177 5148 183
rect 5156 177 5180 183
rect 5197 183 5203 197
rect 5220 197 5276 203
rect 5428 197 5580 203
rect 5844 197 6060 203
rect 6164 197 6204 203
rect 5197 177 5324 183
rect 5364 177 5484 183
rect 5508 177 5644 183
rect 5668 177 5756 183
rect 5789 177 5900 183
rect 4372 157 4403 163
rect 4420 157 4460 163
rect 4484 157 4876 163
rect 5012 157 5052 163
rect 5140 157 5148 163
rect 5204 157 5452 163
rect 5789 163 5795 177
rect 5940 177 5964 183
rect 6180 177 6236 183
rect 5540 157 5795 163
rect 5812 157 6220 163
rect 6260 157 6268 163
rect 3821 144 3827 156
rect 2189 137 2220 143
rect 2324 137 2444 143
rect 2468 137 2492 143
rect 2548 137 3308 143
rect 3316 137 3468 143
rect 3540 137 3580 143
rect 3588 137 3676 143
rect 3684 137 3692 143
rect 3764 137 3820 143
rect 3860 137 4108 143
rect 4132 137 4284 143
rect 4308 137 5036 143
rect 5069 137 5116 143
rect 5069 124 5075 137
rect 5140 137 5308 143
rect 5396 137 5580 143
rect 5716 137 5932 143
rect 5940 137 5996 143
rect 6148 137 6156 143
rect 308 117 380 123
rect 468 117 492 123
rect 820 117 844 123
rect 1172 117 1244 123
rect 1268 117 1276 123
rect 1284 117 1356 123
rect 1460 117 1500 123
rect 1524 117 1564 123
rect 1588 117 1644 123
rect 1668 117 1804 123
rect 1972 117 2028 123
rect 2084 117 2124 123
rect 2148 117 2204 123
rect 2244 117 2476 123
rect 2500 117 2540 123
rect 2548 117 2556 123
rect 2573 117 2620 123
rect 836 97 908 103
rect 916 97 940 103
rect 948 97 1068 103
rect 1076 97 1132 103
rect 1140 97 1228 103
rect 1236 97 1292 103
rect 1316 97 1404 103
rect 1428 97 1852 103
rect 1860 97 1932 103
rect 1956 97 1996 103
rect 2013 97 2060 103
rect 884 77 1020 83
rect 1060 77 1452 83
rect 1469 77 1580 83
rect 1469 63 1475 77
rect 2013 83 2019 97
rect 2100 97 2140 103
rect 2180 97 2268 103
rect 2292 97 2364 103
rect 2573 103 2579 117
rect 2676 117 2899 123
rect 2404 97 2579 103
rect 2596 97 2716 103
rect 2756 97 2812 103
rect 2893 103 2899 117
rect 2916 117 3020 123
rect 3060 117 3507 123
rect 2893 97 3212 103
rect 3236 97 3324 103
rect 3348 97 3372 103
rect 3501 103 3507 117
rect 3524 117 3532 123
rect 3572 117 3676 123
rect 3764 117 3884 123
rect 3892 117 4316 123
rect 4388 117 4396 123
rect 4452 117 4588 123
rect 4596 117 4780 123
rect 4804 117 4812 123
rect 4836 117 4924 123
rect 4948 117 5068 123
rect 5092 117 5180 123
rect 5188 117 5244 123
rect 5332 117 5340 123
rect 5348 117 5388 123
rect 5412 117 5708 123
rect 5748 117 5964 123
rect 6068 117 6092 123
rect 6132 117 6188 123
rect 3501 97 3548 103
rect 3652 97 3852 103
rect 3876 97 3884 103
rect 3908 97 3948 103
rect 3988 97 4044 103
rect 4084 97 4092 103
rect 4116 97 4188 103
rect 4244 97 4492 103
rect 4500 97 5068 103
rect 5076 97 5564 103
rect 5588 97 5628 103
rect 5684 97 5884 103
rect 5908 97 6028 103
rect 2829 84 2835 96
rect 1604 77 2019 83
rect 2036 77 2492 83
rect 2516 77 2540 83
rect 2564 77 2732 83
rect 2756 77 2787 83
rect 580 57 1475 63
rect 1556 57 2140 63
rect 2164 57 2188 63
rect 2212 57 2364 63
rect 2388 57 2764 63
rect 2781 63 2787 77
rect 2852 77 3980 83
rect 4036 77 4044 83
rect 4132 77 4492 83
rect 4516 77 4940 83
rect 4964 77 5196 83
rect 5268 77 5420 83
rect 5476 77 5772 83
rect 5860 77 5932 83
rect 2781 57 2924 63
rect 3092 57 3267 63
rect 244 37 2380 43
rect 2404 37 2556 43
rect 2580 37 2604 43
rect 2628 37 2668 43
rect 2692 37 2828 43
rect 2868 37 2988 43
rect 3044 37 3180 43
rect 3261 43 3267 57
rect 3444 57 3660 63
rect 3684 57 4332 63
rect 4372 57 4412 63
rect 4436 57 4540 63
rect 4564 57 5004 63
rect 5044 57 5212 63
rect 5236 57 5372 63
rect 5460 57 5676 63
rect 5748 57 6028 63
rect 3261 37 3452 43
rect 3476 37 4012 43
rect 4029 37 4188 43
rect 148 17 1548 23
rect 1652 17 2124 23
rect 2148 17 2700 23
rect 2724 17 2828 23
rect 3220 17 3356 23
rect 4029 23 4035 37
rect 4212 37 4668 43
rect 4756 37 5260 43
rect 5284 37 5292 43
rect 5316 37 5788 43
rect 3508 17 4035 23
rect 4148 17 4636 23
rect 4916 17 5356 23
rect 5396 17 5468 23
rect 5492 17 5740 23
rect 5764 17 6124 23
rect 1576 14 1624 16
rect 1576 6 1577 14
rect 1586 6 1587 14
rect 1622 6 1624 14
rect 1576 4 1624 6
rect 4664 14 4712 16
rect 4664 6 4665 14
rect 4674 6 4675 14
rect 4710 6 4712 14
rect 4664 4 4712 6
<< m4contact >>
rect 1708 4616 1716 4624
rect 2412 4616 2420 4624
rect 2732 4616 2740 4624
rect 2892 4616 2900 4624
rect 3020 4616 3028 4624
rect 3244 4616 3252 4624
rect 3308 4616 3316 4624
rect 3468 4616 3476 4624
rect 4460 4616 4468 4624
rect 3114 4606 3121 4614
rect 3121 4606 3122 4614
rect 3126 4606 3131 4614
rect 3131 4606 3133 4614
rect 3133 4606 3134 4614
rect 3138 4606 3141 4614
rect 3141 4606 3143 4614
rect 3143 4606 3146 4614
rect 3150 4606 3151 4614
rect 3151 4606 3158 4614
rect 524 4596 532 4604
rect 2060 4596 2068 4604
rect 2124 4596 2132 4604
rect 2924 4596 2932 4604
rect 748 4576 756 4584
rect 3212 4596 3220 4604
rect 5196 4596 5204 4604
rect 3820 4576 3828 4584
rect 5836 4576 5844 4584
rect 204 4536 212 4544
rect 1132 4536 1140 4544
rect 2540 4556 2548 4564
rect 3628 4556 3636 4564
rect 5596 4556 5604 4564
rect 6156 4556 6164 4564
rect 460 4516 468 4524
rect 716 4516 724 4524
rect 1100 4516 1108 4524
rect 1804 4536 1812 4544
rect 2316 4536 2324 4544
rect 2796 4536 2804 4544
rect 2700 4516 2708 4524
rect 2764 4516 2772 4524
rect 1900 4496 1908 4504
rect 2892 4496 2900 4504
rect 3372 4516 3380 4524
rect 3500 4536 3508 4544
rect 4236 4536 4244 4544
rect 5484 4536 5492 4544
rect 5580 4536 5588 4544
rect 5772 4536 5780 4544
rect 5996 4536 6004 4544
rect 5420 4516 5428 4524
rect 4140 4496 4148 4504
rect 5708 4516 5716 4524
rect 5740 4516 5748 4524
rect 5964 4496 5972 4504
rect 6156 4496 6164 4504
rect 1708 4476 1716 4484
rect 1932 4476 1940 4484
rect 3020 4476 3028 4484
rect 3052 4476 3060 4484
rect 4076 4456 4084 4464
rect 6156 4456 6164 4464
rect 2380 4436 2388 4444
rect 2572 4436 2580 4444
rect 4908 4436 4916 4444
rect 5164 4436 5172 4444
rect 1578 4406 1585 4414
rect 1585 4406 1586 4414
rect 1590 4406 1595 4414
rect 1595 4406 1597 4414
rect 1597 4406 1598 4414
rect 1602 4406 1605 4414
rect 1605 4406 1607 4414
rect 1607 4406 1610 4414
rect 1614 4406 1615 4414
rect 1615 4406 1622 4414
rect 4666 4406 4673 4414
rect 4673 4406 4674 4414
rect 4678 4406 4683 4414
rect 4683 4406 4685 4414
rect 4685 4406 4686 4414
rect 4690 4406 4693 4414
rect 4693 4406 4695 4414
rect 4695 4406 4698 4414
rect 4702 4406 4703 4414
rect 4703 4406 4710 4414
rect 1772 4396 1780 4404
rect 3788 4396 3796 4404
rect 1260 4376 1268 4384
rect 236 4356 244 4364
rect 1516 4356 1524 4364
rect 1932 4376 1940 4384
rect 2956 4376 2964 4384
rect 5356 4376 5364 4384
rect 5388 4376 5396 4384
rect 2316 4356 2324 4364
rect 2796 4356 2804 4364
rect 3596 4356 3604 4364
rect 1740 4336 1748 4344
rect 3404 4336 3412 4344
rect 3500 4336 3508 4344
rect 3692 4336 3700 4344
rect 5516 4336 5524 4344
rect 6252 4336 6260 4344
rect 1004 4316 1012 4324
rect 2444 4316 2452 4324
rect 4204 4316 4212 4324
rect 5484 4316 5492 4324
rect 5580 4316 5588 4324
rect 1772 4296 1780 4304
rect 2860 4296 2868 4304
rect 3020 4296 3028 4304
rect 3436 4296 3444 4304
rect 3564 4296 3572 4304
rect 4268 4296 4276 4304
rect 4300 4296 4308 4304
rect 4492 4296 4500 4304
rect 5900 4296 5908 4304
rect 1964 4276 1972 4284
rect 1996 4276 2004 4284
rect 2028 4276 2036 4284
rect 2188 4276 2196 4284
rect 2332 4276 2340 4284
rect 1036 4256 1044 4264
rect 1420 4256 1428 4264
rect 3724 4276 3732 4284
rect 4076 4276 4084 4284
rect 5420 4276 5428 4284
rect 5484 4276 5492 4284
rect 2924 4256 2932 4264
rect 2988 4256 2996 4264
rect 3500 4256 3508 4264
rect 3596 4256 3604 4264
rect 5932 4256 5940 4264
rect 6028 4256 6036 4264
rect 6124 4256 6132 4264
rect 812 4236 820 4244
rect 876 4236 884 4244
rect 1708 4236 1716 4244
rect 2508 4236 2516 4244
rect 3628 4236 3636 4244
rect 5388 4236 5396 4244
rect 5676 4236 5684 4244
rect 1388 4216 1396 4224
rect 2092 4216 2100 4224
rect 2412 4216 2420 4224
rect 2924 4216 2932 4224
rect 3308 4216 3316 4224
rect 3404 4216 3412 4224
rect 3980 4216 3988 4224
rect 4588 4216 4596 4224
rect 3114 4206 3121 4214
rect 3121 4206 3122 4214
rect 3126 4206 3131 4214
rect 3131 4206 3133 4214
rect 3133 4206 3134 4214
rect 3138 4206 3141 4214
rect 3141 4206 3143 4214
rect 3143 4206 3146 4214
rect 3150 4206 3151 4214
rect 3151 4206 3158 4214
rect 364 4176 372 4184
rect 364 4156 372 4164
rect 972 4176 980 4184
rect 2028 4176 2036 4184
rect 2348 4176 2356 4184
rect 2380 4176 2388 4184
rect 876 4156 884 4164
rect 1660 4156 1668 4164
rect 4076 4196 4084 4204
rect 4012 4176 4020 4184
rect 4204 4176 4212 4184
rect 4396 4196 4404 4204
rect 5420 4196 5428 4204
rect 5868 4216 5876 4224
rect 5676 4176 5684 4184
rect 2636 4156 2644 4164
rect 3340 4156 3348 4164
rect 3692 4156 3700 4164
rect 684 4136 692 4144
rect 1036 4136 1044 4144
rect 1356 4136 1364 4144
rect 140 4116 148 4124
rect 204 4116 212 4124
rect 204 4096 212 4104
rect 332 4096 340 4104
rect 1228 4116 1236 4124
rect 1260 4116 1268 4124
rect 1420 4136 1428 4144
rect 2060 4116 2068 4124
rect 2412 4116 2420 4124
rect 2444 4116 2452 4124
rect 2668 4116 2676 4124
rect 3404 4136 3412 4144
rect 4364 4156 4372 4164
rect 5036 4156 5044 4164
rect 5260 4156 5268 4164
rect 5932 4156 5940 4164
rect 6124 4156 6132 4164
rect 6188 4156 6196 4164
rect 3020 4116 3028 4124
rect 3340 4116 3348 4124
rect 3980 4116 3988 4124
rect 4204 4136 4212 4144
rect 4236 4136 4244 4144
rect 4300 4136 4308 4144
rect 5676 4136 5684 4144
rect 5292 4116 5300 4124
rect 5708 4116 5716 4124
rect 5836 4116 5844 4124
rect 6220 4116 6228 4124
rect 1004 4096 1012 4104
rect 1676 4096 1684 4104
rect 1964 4096 1972 4104
rect 2188 4096 2196 4104
rect 2380 4096 2388 4104
rect 2508 4096 2516 4104
rect 3308 4096 3316 4104
rect 4396 4096 4404 4104
rect 5164 4096 5172 4104
rect 5740 4096 5748 4104
rect 460 4076 468 4084
rect 1836 4076 1844 4084
rect 1868 4076 1876 4084
rect 2412 4076 2420 4084
rect 2572 4076 2580 4084
rect 2892 4076 2900 4084
rect 3276 4076 3284 4084
rect 3660 4076 3668 4084
rect 3980 4076 3988 4084
rect 4300 4076 4308 4084
rect 5868 4076 5876 4084
rect 6028 4076 6036 4084
rect 6092 4076 6100 4084
rect 6284 4076 6292 4084
rect 1228 4056 1236 4064
rect 1324 4056 1332 4064
rect 1356 4056 1364 4064
rect 1804 4056 1812 4064
rect 1932 4056 1940 4064
rect 1292 4036 1300 4044
rect 1516 4036 1524 4044
rect 1708 4036 1716 4044
rect 1820 4036 1828 4044
rect 1996 4056 2004 4064
rect 2988 4056 2996 4064
rect 4236 4056 4244 4064
rect 4268 4056 4276 4064
rect 4556 4056 4564 4064
rect 5836 4056 5844 4064
rect 2316 4036 2324 4044
rect 2380 4036 2388 4044
rect 2572 4036 2580 4044
rect 1228 4016 1236 4024
rect 1484 4016 1492 4024
rect 2028 4016 2036 4024
rect 2156 4016 2164 4024
rect 2636 4016 2644 4024
rect 2828 4016 2836 4024
rect 4620 4016 4628 4024
rect 5228 4016 5236 4024
rect 5356 4016 5364 4024
rect 6124 4036 6132 4044
rect 1578 4006 1585 4014
rect 1585 4006 1586 4014
rect 1590 4006 1595 4014
rect 1595 4006 1597 4014
rect 1597 4006 1598 4014
rect 1602 4006 1605 4014
rect 1605 4006 1607 4014
rect 1607 4006 1610 4014
rect 1614 4006 1615 4014
rect 1615 4006 1622 4014
rect 4666 4006 4673 4014
rect 4673 4006 4674 4014
rect 4678 4006 4683 4014
rect 4683 4006 4685 4014
rect 4685 4006 4686 4014
rect 4690 4006 4693 4014
rect 4693 4006 4695 4014
rect 4695 4006 4698 4014
rect 4702 4006 4703 4014
rect 4703 4006 4710 4014
rect 1516 3996 1524 4004
rect 2732 3996 2740 4004
rect 2860 3996 2868 4004
rect 3532 3996 3540 4004
rect 3660 3996 3668 4004
rect 3692 3996 3700 4004
rect 3884 3996 3892 4004
rect 4012 3996 4020 4004
rect 4172 3996 4180 4004
rect 4428 3996 4436 4004
rect 4460 3996 4468 4004
rect 1196 3976 1204 3984
rect 1388 3976 1396 3984
rect 1452 3976 1460 3984
rect 1132 3956 1140 3964
rect 1164 3956 1172 3964
rect 1868 3976 1876 3984
rect 2060 3976 2068 3984
rect 2444 3976 2452 3984
rect 2604 3976 2612 3984
rect 2764 3976 2772 3984
rect 2796 3976 2804 3984
rect 3372 3976 3380 3984
rect 4140 3976 4148 3984
rect 4588 3976 4596 3984
rect 4780 3976 4788 3984
rect 6060 3976 6068 3984
rect 2476 3956 2484 3964
rect 2860 3956 2868 3964
rect 3564 3956 3572 3964
rect 3948 3956 3956 3964
rect 4364 3956 4372 3964
rect 1452 3936 1460 3944
rect 2028 3936 2036 3944
rect 2444 3936 2452 3944
rect 2636 3936 2644 3944
rect 2700 3936 2708 3944
rect 3436 3940 3444 3948
rect 3596 3936 3604 3944
rect 4012 3936 4020 3944
rect 4076 3936 4084 3944
rect 4140 3936 4148 3944
rect 5388 3936 5396 3944
rect 5932 3936 5940 3944
rect 204 3916 212 3924
rect 172 3896 180 3904
rect 236 3876 244 3884
rect 332 3916 340 3924
rect 524 3916 532 3924
rect 1260 3916 1268 3924
rect 1484 3916 1492 3924
rect 1868 3916 1876 3924
rect 1996 3916 2004 3924
rect 2156 3916 2164 3924
rect 2540 3916 2548 3924
rect 2732 3916 2740 3924
rect 2764 3916 2772 3924
rect 2860 3916 2868 3924
rect 3340 3916 3348 3924
rect 3404 3916 3412 3924
rect 3436 3912 3444 3920
rect 3980 3916 3988 3924
rect 4108 3916 4116 3924
rect 4172 3916 4180 3924
rect 4460 3916 4468 3924
rect 5228 3916 5236 3924
rect 5580 3916 5588 3924
rect 6156 3916 6164 3924
rect 556 3896 564 3904
rect 524 3876 532 3884
rect 140 3856 148 3864
rect 204 3856 212 3864
rect 972 3856 980 3864
rect 1068 3856 1076 3864
rect 1196 3856 1204 3864
rect 1548 3876 1556 3884
rect 2060 3896 2068 3904
rect 2316 3896 2324 3904
rect 2380 3896 2388 3904
rect 2988 3896 2996 3904
rect 3212 3896 3220 3904
rect 3308 3896 3316 3904
rect 3500 3896 3508 3904
rect 3660 3896 3668 3904
rect 3756 3896 3764 3904
rect 3852 3896 3860 3904
rect 1804 3876 1812 3884
rect 1836 3876 1844 3884
rect 2572 3876 2580 3884
rect 2668 3876 2676 3884
rect 2796 3876 2804 3884
rect 3564 3876 3572 3884
rect 3692 3876 3700 3884
rect 3724 3876 3732 3884
rect 5260 3896 5268 3904
rect 5740 3896 5748 3904
rect 5772 3896 5780 3904
rect 6124 3896 6132 3904
rect 5228 3876 5236 3884
rect 6188 3876 6196 3884
rect 1004 3836 1012 3844
rect 1228 3836 1236 3844
rect 1260 3836 1268 3844
rect 1516 3856 1524 3864
rect 1804 3836 1812 3844
rect 2892 3856 2900 3864
rect 3756 3856 3764 3864
rect 4140 3856 4148 3864
rect 5356 3856 5364 3864
rect 5708 3856 5716 3864
rect 2060 3836 2068 3844
rect 812 3816 820 3824
rect 3212 3836 3220 3844
rect 3244 3836 3252 3844
rect 3308 3836 3316 3844
rect 3340 3836 3348 3844
rect 3628 3836 3636 3844
rect 3692 3836 3700 3844
rect 3852 3836 3860 3844
rect 6028 3836 6036 3844
rect 3404 3816 3412 3824
rect 5292 3816 5300 3824
rect 5836 3816 5844 3824
rect 6156 3816 6164 3824
rect 3114 3806 3121 3814
rect 3121 3806 3122 3814
rect 3126 3806 3131 3814
rect 3131 3806 3133 3814
rect 3133 3806 3134 3814
rect 3138 3806 3141 3814
rect 3141 3806 3143 3814
rect 3143 3806 3146 3814
rect 3150 3806 3151 3814
rect 3151 3806 3158 3814
rect 268 3796 276 3804
rect 396 3796 404 3804
rect 476 3796 484 3804
rect 940 3796 948 3804
rect 1420 3796 1428 3804
rect 1708 3796 1716 3804
rect 1740 3796 1748 3804
rect 1772 3780 1780 3788
rect 2220 3796 2228 3804
rect 3052 3796 3060 3804
rect 4172 3796 4180 3804
rect 5452 3796 5460 3804
rect 6188 3796 6196 3804
rect 2508 3776 2516 3784
rect 2540 3776 2548 3784
rect 4268 3776 4276 3784
rect 5676 3776 5684 3784
rect 5804 3776 5812 3784
rect 5836 3776 5844 3784
rect 6060 3776 6068 3784
rect 6124 3776 6132 3784
rect 300 3756 308 3764
rect 908 3756 916 3764
rect 1132 3756 1140 3764
rect 1196 3756 1204 3764
rect 1420 3756 1428 3764
rect 1772 3752 1780 3760
rect 1900 3756 1908 3764
rect 2924 3756 2932 3764
rect 3180 3756 3188 3764
rect 3468 3756 3476 3764
rect 3532 3756 3540 3764
rect 140 3736 148 3744
rect 204 3736 212 3744
rect 396 3736 404 3744
rect 460 3736 468 3744
rect 364 3716 372 3724
rect 620 3716 628 3724
rect 1388 3716 1396 3724
rect 204 3696 212 3704
rect 236 3696 244 3704
rect 556 3696 564 3704
rect 1132 3696 1140 3704
rect 2444 3736 2452 3744
rect 1452 3716 1460 3724
rect 1548 3716 1556 3724
rect 1484 3696 1492 3704
rect 1676 3696 1684 3704
rect 1740 3696 1748 3704
rect 1804 3716 1812 3724
rect 2316 3716 2324 3724
rect 2764 3716 2772 3724
rect 2860 3716 2868 3724
rect 3628 3736 3636 3744
rect 3276 3716 3284 3724
rect 3820 3756 3828 3764
rect 4012 3756 4020 3764
rect 4908 3756 4916 3764
rect 5484 3756 5492 3764
rect 5548 3756 5556 3764
rect 5900 3756 5908 3764
rect 5932 3756 5940 3764
rect 4108 3736 4116 3744
rect 2092 3696 2100 3704
rect 2188 3696 2196 3704
rect 2284 3696 2292 3704
rect 2604 3696 2612 3704
rect 2732 3696 2740 3704
rect 2828 3696 2836 3704
rect 3020 3696 3028 3704
rect 2252 3676 2260 3684
rect 2380 3676 2388 3684
rect 2444 3676 2452 3684
rect 2508 3676 2516 3684
rect 3628 3696 3636 3704
rect 3788 3716 3796 3724
rect 4044 3716 4052 3724
rect 5324 3736 5332 3744
rect 5644 3736 5652 3744
rect 6284 3756 6292 3764
rect 4236 3716 4244 3724
rect 4556 3716 4564 3724
rect 4588 3716 4596 3724
rect 5740 3716 5748 3724
rect 6156 3716 6164 3724
rect 3980 3696 3988 3704
rect 4012 3696 4020 3704
rect 5292 3696 5300 3704
rect 5324 3696 5332 3704
rect 5708 3696 5716 3704
rect 5836 3696 5844 3704
rect 6028 3696 6036 3704
rect 6284 3696 6292 3704
rect 3244 3676 3252 3684
rect 428 3656 436 3664
rect 460 3656 468 3664
rect 1036 3656 1044 3664
rect 2348 3656 2356 3664
rect 2764 3656 2772 3664
rect 2860 3656 2868 3664
rect 3276 3656 3284 3664
rect 3436 3656 3444 3664
rect 3852 3676 3860 3684
rect 4076 3676 4084 3684
rect 4396 3676 4404 3684
rect 4620 3676 4628 3684
rect 5612 3676 5620 3684
rect 6124 3676 6132 3684
rect 140 3636 148 3644
rect 972 3636 980 3644
rect 1836 3636 1844 3644
rect 2604 3636 2612 3644
rect 5324 3636 5332 3644
rect 236 3616 244 3624
rect 1388 3616 1396 3624
rect 1676 3616 1684 3624
rect 2028 3616 2036 3624
rect 2668 3616 2676 3624
rect 3180 3616 3188 3624
rect 3436 3616 3444 3624
rect 3660 3616 3668 3624
rect 4172 3616 4180 3624
rect 4236 3616 4244 3624
rect 5228 3616 5236 3624
rect 5580 3616 5588 3624
rect 5836 3616 5844 3624
rect 1578 3606 1585 3614
rect 1585 3606 1586 3614
rect 1590 3606 1595 3614
rect 1595 3606 1597 3614
rect 1597 3606 1598 3614
rect 1602 3606 1605 3614
rect 1605 3606 1607 3614
rect 1607 3606 1610 3614
rect 1614 3606 1615 3614
rect 1615 3606 1622 3614
rect 4666 3606 4673 3614
rect 4673 3606 4674 3614
rect 4678 3606 4683 3614
rect 4683 3606 4685 3614
rect 4685 3606 4686 3614
rect 4690 3606 4693 3614
rect 4693 3606 4695 3614
rect 4695 3606 4698 3614
rect 4702 3606 4703 3614
rect 4703 3606 4710 3614
rect 140 3596 148 3604
rect 812 3576 820 3584
rect 1132 3596 1140 3604
rect 1164 3576 1172 3584
rect 1836 3596 1844 3604
rect 1868 3596 1876 3604
rect 2508 3596 2516 3604
rect 2572 3596 2580 3604
rect 2764 3596 2772 3604
rect 2860 3596 2868 3604
rect 2908 3596 2916 3604
rect 3052 3596 3060 3604
rect 3820 3596 3828 3604
rect 4044 3596 4052 3604
rect 6092 3596 6100 3604
rect 2220 3576 2228 3584
rect 2412 3576 2420 3584
rect 844 3556 852 3564
rect 1196 3556 1204 3564
rect 268 3536 276 3544
rect 556 3536 564 3544
rect 1484 3536 1492 3544
rect 1548 3536 1556 3544
rect 204 3516 212 3524
rect 396 3516 404 3524
rect 588 3516 596 3524
rect 652 3516 660 3524
rect 908 3516 916 3524
rect 1260 3516 1268 3524
rect 1324 3516 1332 3524
rect 1356 3516 1364 3524
rect 1388 3516 1396 3524
rect 1420 3516 1428 3524
rect 1708 3556 1716 3564
rect 1900 3556 1908 3564
rect 2028 3556 2036 3564
rect 2444 3556 2452 3564
rect 2540 3556 2548 3564
rect 2732 3556 2740 3564
rect 3212 3556 3220 3564
rect 3756 3556 3764 3564
rect 3820 3556 3828 3564
rect 4012 3556 4020 3564
rect 1964 3536 1972 3544
rect 1996 3536 2004 3544
rect 2316 3536 2324 3544
rect 3308 3536 3316 3544
rect 4172 3536 4180 3544
rect 5228 3536 5236 3544
rect 268 3496 276 3504
rect 1516 3496 1524 3504
rect 620 3476 628 3484
rect 1356 3476 1364 3484
rect 1484 3476 1492 3484
rect 1804 3496 1812 3504
rect 2348 3516 2356 3524
rect 1708 3476 1716 3484
rect 1772 3476 1780 3484
rect 1868 3476 1876 3484
rect 2188 3496 2196 3504
rect 2412 3496 2420 3504
rect 2476 3496 2484 3504
rect 2940 3516 2948 3524
rect 2988 3516 2996 3524
rect 3980 3516 3988 3524
rect 4460 3516 4468 3524
rect 5420 3516 5428 3524
rect 5484 3516 5492 3524
rect 5772 3536 5780 3544
rect 5868 3536 5876 3544
rect 5964 3536 5972 3544
rect 5804 3516 5812 3524
rect 5836 3516 5844 3524
rect 716 3456 724 3464
rect 1164 3456 1172 3464
rect 1964 3456 1972 3464
rect 2220 3476 2228 3484
rect 2252 3476 2260 3484
rect 2636 3476 2644 3484
rect 3340 3496 3348 3504
rect 3628 3496 3636 3504
rect 3852 3496 3860 3504
rect 3948 3496 3956 3504
rect 4780 3496 4788 3504
rect 5932 3496 5940 3504
rect 2988 3476 2996 3484
rect 3036 3476 3044 3484
rect 2092 3436 2100 3444
rect 2700 3456 2708 3464
rect 3308 3456 3316 3464
rect 1260 3416 1268 3424
rect 2316 3416 2324 3424
rect 3468 3476 3476 3484
rect 3660 3476 3668 3484
rect 3756 3476 3764 3484
rect 4268 3476 4276 3484
rect 5612 3476 5620 3484
rect 5708 3476 5716 3484
rect 5964 3476 5972 3484
rect 3564 3456 3572 3464
rect 3788 3456 3796 3464
rect 4588 3456 4596 3464
rect 5420 3456 5428 3464
rect 5740 3456 5748 3464
rect 6124 3456 6132 3464
rect 3756 3436 3764 3444
rect 3916 3436 3924 3444
rect 3948 3436 3956 3444
rect 5676 3436 5684 3444
rect 5964 3436 5972 3444
rect 6092 3436 6100 3444
rect 492 3396 500 3404
rect 940 3396 948 3404
rect 1100 3396 1108 3404
rect 1196 3396 1204 3404
rect 1324 3396 1332 3404
rect 1836 3396 1844 3404
rect 1964 3396 1972 3404
rect 2092 3396 2100 3404
rect 2412 3396 2420 3404
rect 2924 3416 2932 3424
rect 2956 3416 2964 3424
rect 3596 3416 3604 3424
rect 3628 3416 3636 3424
rect 3114 3406 3121 3414
rect 3121 3406 3122 3414
rect 3126 3406 3131 3414
rect 3131 3406 3133 3414
rect 3133 3406 3134 3414
rect 3138 3406 3141 3414
rect 3141 3406 3143 3414
rect 3143 3406 3146 3414
rect 3150 3406 3151 3414
rect 3151 3406 3158 3414
rect 2476 3396 2484 3404
rect 524 3376 532 3384
rect 876 3376 884 3384
rect 1132 3376 1140 3384
rect 1228 3376 1236 3384
rect 1260 3376 1268 3384
rect 1420 3376 1428 3384
rect 2636 3376 2644 3384
rect 2924 3376 2932 3384
rect 2956 3376 2964 3384
rect 3244 3396 3252 3404
rect 3628 3396 3636 3404
rect 5836 3416 5844 3424
rect 5580 3396 5588 3404
rect 5740 3396 5748 3404
rect 5964 3396 5972 3404
rect 3276 3376 3284 3384
rect 3372 3376 3380 3384
rect 3500 3376 3508 3384
rect 5356 3376 5364 3384
rect 5548 3376 5556 3384
rect 6188 3376 6196 3384
rect 588 3356 596 3364
rect 844 3356 852 3364
rect 1324 3356 1332 3364
rect 1900 3356 1908 3364
rect 1996 3356 2004 3364
rect 908 3336 916 3344
rect 1004 3336 1012 3344
rect 1036 3336 1044 3344
rect 2316 3356 2324 3364
rect 2252 3336 2260 3344
rect 2380 3336 2388 3344
rect 2412 3336 2420 3344
rect 2572 3356 2580 3364
rect 2988 3356 2996 3364
rect 3084 3356 3092 3364
rect 3244 3356 3252 3364
rect 3692 3356 3700 3364
rect 3756 3356 3764 3364
rect 5452 3356 5460 3364
rect 6124 3356 6132 3364
rect 620 3316 628 3324
rect 556 3276 564 3284
rect 1164 3316 1172 3324
rect 1516 3316 1524 3324
rect 1676 3316 1684 3324
rect 1708 3316 1716 3324
rect 1804 3316 1812 3324
rect 1836 3316 1844 3324
rect 2124 3316 2132 3324
rect 2540 3316 2548 3324
rect 2956 3336 2964 3344
rect 3212 3336 3220 3344
rect 3468 3336 3476 3344
rect 3532 3336 3540 3344
rect 3820 3336 3828 3344
rect 3884 3336 3892 3344
rect 5164 3336 5172 3344
rect 5644 3336 5652 3344
rect 6188 3336 6196 3344
rect 2668 3316 2676 3324
rect 3372 3316 3380 3324
rect 3404 3316 3412 3324
rect 3628 3316 3636 3324
rect 3852 3316 3860 3324
rect 3916 3316 3924 3324
rect 4492 3316 4500 3324
rect 1388 3296 1396 3304
rect 1932 3296 1940 3304
rect 1964 3296 1972 3304
rect 2060 3296 2068 3304
rect 3052 3296 3060 3304
rect 3084 3296 3092 3304
rect 3180 3296 3188 3304
rect 4268 3296 4276 3304
rect 5164 3296 5172 3304
rect 5324 3296 5332 3304
rect 5516 3316 5524 3324
rect 5900 3316 5908 3324
rect 6156 3296 6164 3304
rect 6188 3296 6196 3304
rect 1548 3276 1556 3284
rect 5260 3276 5268 3284
rect 6124 3276 6132 3284
rect 812 3256 820 3264
rect 1708 3256 1716 3264
rect 1740 3256 1748 3264
rect 1772 3256 1780 3264
rect 2028 3256 2036 3264
rect 2156 3256 2164 3264
rect 2348 3256 2356 3264
rect 2732 3256 2740 3264
rect 2860 3256 2868 3264
rect 2924 3256 2932 3264
rect 12 3236 20 3244
rect 268 3216 276 3224
rect 428 3216 436 3224
rect 1004 3236 1012 3244
rect 1068 3236 1076 3244
rect 1900 3236 1908 3244
rect 2092 3236 2100 3244
rect 2124 3236 2132 3244
rect 2828 3236 2836 3244
rect 3084 3236 3092 3244
rect 5356 3256 5364 3264
rect 5388 3256 5396 3264
rect 3420 3236 3428 3244
rect 3852 3236 3860 3244
rect 5580 3236 5588 3244
rect 1196 3216 1204 3224
rect 1516 3216 1524 3224
rect 1772 3216 1780 3224
rect 2284 3216 2292 3224
rect 2508 3216 2516 3224
rect 1578 3206 1585 3214
rect 1585 3206 1586 3214
rect 1590 3206 1595 3214
rect 1595 3206 1597 3214
rect 1597 3206 1598 3214
rect 1602 3206 1605 3214
rect 1605 3206 1607 3214
rect 1607 3206 1610 3214
rect 1614 3206 1615 3214
rect 1615 3206 1622 3214
rect 140 3196 148 3204
rect 1228 3196 1236 3204
rect 1260 3196 1268 3204
rect 1420 3196 1428 3204
rect 2220 3196 2228 3204
rect 2860 3216 2868 3224
rect 2956 3216 2964 3224
rect 3372 3216 3380 3224
rect 3404 3216 3412 3224
rect 4108 3216 4116 3224
rect 4236 3216 4244 3224
rect 4666 3206 4673 3214
rect 4673 3206 4674 3214
rect 4678 3206 4683 3214
rect 4683 3206 4685 3214
rect 4685 3206 4686 3214
rect 4690 3206 4693 3214
rect 4693 3206 4695 3214
rect 4695 3206 4698 3214
rect 4702 3206 4703 3214
rect 4703 3206 4710 3214
rect 2572 3196 2580 3204
rect 3980 3196 3988 3204
rect 4012 3196 4020 3204
rect 5388 3196 5396 3204
rect 844 3176 852 3184
rect 1036 3176 1044 3184
rect 1068 3176 1076 3184
rect 1292 3176 1300 3184
rect 140 3156 148 3164
rect 556 3136 564 3144
rect 588 3156 596 3164
rect 940 3156 948 3164
rect 1212 3156 1220 3164
rect 1324 3156 1332 3164
rect 2092 3176 2100 3184
rect 2796 3176 2804 3184
rect 3244 3176 3252 3184
rect 3436 3176 3444 3184
rect 3468 3176 3476 3184
rect 4332 3176 4340 3184
rect 5196 3176 5204 3184
rect 5804 3176 5812 3184
rect 1292 3136 1300 3144
rect 460 3116 468 3124
rect 588 3116 596 3124
rect 1196 3116 1204 3124
rect 1244 3116 1252 3124
rect 1420 3116 1428 3124
rect 1644 3136 1652 3144
rect 1676 3116 1684 3124
rect 2060 3136 2068 3144
rect 2444 3156 2452 3164
rect 2508 3156 2516 3164
rect 2636 3156 2644 3164
rect 2668 3156 2676 3164
rect 2732 3156 2740 3164
rect 3404 3156 3412 3164
rect 3692 3156 3700 3164
rect 3820 3156 3828 3164
rect 4140 3156 4148 3164
rect 5932 3156 5940 3164
rect 2956 3136 2964 3144
rect 4044 3136 4052 3144
rect 5548 3136 5556 3144
rect 236 3096 244 3104
rect 332 3096 340 3104
rect 620 3096 628 3104
rect 908 3096 916 3104
rect 972 3096 980 3104
rect 1036 3096 1044 3104
rect 204 3076 212 3084
rect 588 3076 596 3084
rect 876 3076 884 3084
rect 1260 3096 1268 3104
rect 1484 3096 1492 3104
rect 1772 3096 1780 3104
rect 1836 3096 1844 3104
rect 2124 3096 2132 3104
rect 2156 3096 2164 3104
rect 2444 3116 2452 3124
rect 3084 3116 3092 3124
rect 3724 3116 3732 3124
rect 3916 3116 3924 3124
rect 4172 3116 4180 3124
rect 6188 3116 6196 3124
rect 2476 3096 2484 3104
rect 2636 3096 2644 3104
rect 2796 3096 2804 3104
rect 2828 3096 2836 3104
rect 1196 3076 1204 3084
rect 1388 3076 1396 3084
rect 780 3056 788 3064
rect 972 3056 980 3064
rect 1324 3056 1332 3064
rect 1532 3076 1540 3084
rect 1740 3076 1748 3084
rect 1804 3076 1812 3084
rect 2380 3076 2388 3084
rect 2508 3076 2516 3084
rect 2604 3076 2612 3084
rect 2636 3076 2644 3084
rect 1356 3036 1364 3044
rect 492 3016 500 3024
rect 844 3016 852 3024
rect 1708 3056 1716 3064
rect 1836 3056 1844 3064
rect 1900 3056 1908 3064
rect 1996 3056 2004 3064
rect 2028 3056 2036 3064
rect 2348 3056 2356 3064
rect 2444 3056 2452 3064
rect 2732 3076 2740 3084
rect 2988 3076 2996 3084
rect 3020 3076 3028 3084
rect 3532 3096 3540 3104
rect 3276 3076 3284 3084
rect 3340 3076 3348 3084
rect 5644 3096 5652 3104
rect 5932 3096 5940 3104
rect 3660 3076 3668 3084
rect 3708 3076 3716 3084
rect 3788 3076 3796 3084
rect 3884 3076 3892 3084
rect 3180 3056 3188 3064
rect 2156 3036 2164 3044
rect 2540 3036 2548 3044
rect 2636 3036 2644 3044
rect 1676 3016 1684 3024
rect 1900 3016 1908 3024
rect 1932 3016 1940 3024
rect 2188 3016 2196 3024
rect 2284 3016 2292 3024
rect 2508 3016 2516 3024
rect 2796 3016 2804 3024
rect 3020 3036 3028 3044
rect 3244 3036 3252 3044
rect 3404 3056 3412 3064
rect 3372 3036 3380 3044
rect 3596 3056 3604 3064
rect 4060 3076 4068 3084
rect 4300 3076 4308 3084
rect 5164 3076 5172 3084
rect 5676 3076 5684 3084
rect 5900 3076 5908 3084
rect 3980 3056 3988 3064
rect 3500 3036 3508 3044
rect 4204 3036 4212 3044
rect 4524 3036 4532 3044
rect 5196 3056 5204 3064
rect 5324 3056 5332 3064
rect 5420 3056 5428 3064
rect 5484 3056 5492 3064
rect 5644 3056 5652 3064
rect 3308 3016 3316 3024
rect 4140 3016 4148 3024
rect 4428 3016 4436 3024
rect 5388 3016 5396 3024
rect 5548 3016 5556 3024
rect 6124 3016 6132 3024
rect 3114 3006 3121 3014
rect 3121 3006 3122 3014
rect 3126 3006 3131 3014
rect 3131 3006 3133 3014
rect 3133 3006 3134 3014
rect 3138 3006 3141 3014
rect 3141 3006 3143 3014
rect 3143 3006 3146 3014
rect 3150 3006 3151 3014
rect 3151 3006 3158 3014
rect 588 2996 596 3004
rect 716 2996 724 3004
rect 1452 2996 1460 3004
rect 1516 2996 1524 3004
rect 1644 2996 1652 3004
rect 1868 2996 1876 3004
rect 2156 2996 2164 3004
rect 2540 2996 2548 3004
rect 2604 2996 2612 3004
rect 2732 2996 2740 3004
rect 2892 2996 2900 3004
rect 2924 2996 2932 3004
rect 2956 2996 2964 3004
rect 2988 2996 2996 3004
rect 3340 2996 3348 3004
rect 3404 2996 3412 3004
rect 3436 2996 3444 3004
rect 3660 2996 3668 3004
rect 3692 2996 3700 3004
rect 4012 2996 4020 3004
rect 4076 2996 4084 3004
rect 5228 2996 5236 3004
rect 684 2976 692 2984
rect 1228 2976 1236 2984
rect 1420 2976 1428 2984
rect 1452 2976 1460 2984
rect 3852 2976 3860 2984
rect 5804 2976 5812 2984
rect 332 2956 340 2964
rect 780 2956 788 2964
rect 1164 2956 1172 2964
rect 876 2936 884 2944
rect 1004 2936 1012 2944
rect 1068 2936 1076 2944
rect 1324 2936 1332 2944
rect 1804 2956 1812 2964
rect 1996 2956 2004 2964
rect 2476 2956 2484 2964
rect 2668 2956 2676 2964
rect 2732 2956 2740 2964
rect 2796 2956 2804 2964
rect 1420 2936 1428 2944
rect 2188 2936 2196 2944
rect 2220 2936 2228 2944
rect 2444 2936 2452 2944
rect 2764 2936 2772 2944
rect 3084 2956 3092 2964
rect 3404 2956 3412 2964
rect 3468 2956 3476 2964
rect 3276 2936 3284 2944
rect 3308 2936 3316 2944
rect 3372 2936 3380 2944
rect 4044 2956 4052 2964
rect 3724 2936 3732 2944
rect 4364 2956 4372 2964
rect 5228 2956 5236 2964
rect 5484 2956 5492 2964
rect 6188 2956 6196 2964
rect 4236 2936 4244 2944
rect 5292 2936 5300 2944
rect 5644 2936 5652 2944
rect 5804 2936 5812 2944
rect 396 2916 404 2924
rect 492 2916 500 2924
rect 1036 2916 1044 2924
rect 1132 2916 1140 2924
rect 908 2896 916 2904
rect 1164 2896 1172 2904
rect 1260 2916 1268 2924
rect 460 2876 468 2884
rect 1068 2876 1076 2884
rect 1484 2896 1492 2904
rect 1548 2896 1556 2904
rect 1740 2916 1748 2924
rect 1836 2896 1844 2904
rect 1868 2876 1876 2884
rect 2092 2876 2100 2884
rect 2284 2896 2292 2904
rect 2348 2876 2356 2884
rect 2732 2916 2740 2924
rect 2668 2896 2676 2904
rect 3420 2916 3428 2924
rect 3724 2916 3732 2924
rect 3916 2916 3924 2924
rect 3948 2916 3956 2924
rect 4364 2916 4372 2924
rect 4588 2916 4596 2924
rect 5260 2916 5268 2924
rect 5612 2916 5620 2924
rect 2764 2876 2772 2884
rect 3276 2896 3284 2904
rect 3532 2896 3540 2904
rect 4300 2896 4308 2904
rect 5164 2896 5172 2904
rect 5740 2916 5748 2924
rect 6188 2896 6196 2904
rect 2988 2876 2996 2884
rect 3052 2876 3060 2884
rect 3660 2876 3668 2884
rect 5804 2876 5812 2884
rect 1740 2856 1748 2864
rect 1804 2856 1812 2864
rect 2252 2856 2260 2864
rect 2540 2856 2548 2864
rect 2636 2856 2644 2864
rect 1228 2836 1236 2844
rect 1292 2836 1300 2844
rect 1772 2836 1780 2844
rect 1868 2836 1876 2844
rect 2700 2836 2708 2844
rect 2892 2836 2900 2844
rect 3468 2856 3476 2864
rect 3596 2856 3604 2864
rect 4140 2856 4148 2864
rect 5228 2856 5236 2864
rect 5324 2856 5332 2864
rect 3244 2836 3252 2844
rect 3404 2836 3412 2844
rect 3436 2836 3444 2844
rect 236 2816 244 2824
rect 652 2816 660 2824
rect 844 2816 852 2824
rect 1260 2816 1268 2824
rect 1964 2816 1972 2824
rect 2444 2816 2452 2824
rect 2860 2816 2868 2824
rect 5772 2836 5780 2844
rect 4620 2816 4628 2824
rect 5804 2816 5812 2824
rect 1578 2806 1585 2814
rect 1585 2806 1586 2814
rect 1590 2806 1595 2814
rect 1595 2806 1597 2814
rect 1597 2806 1598 2814
rect 1602 2806 1605 2814
rect 1605 2806 1607 2814
rect 1607 2806 1610 2814
rect 1614 2806 1615 2814
rect 1615 2806 1622 2814
rect 4666 2806 4673 2814
rect 4673 2806 4674 2814
rect 4678 2806 4683 2814
rect 4683 2806 4685 2814
rect 4685 2806 4686 2814
rect 4690 2806 4693 2814
rect 4693 2806 4695 2814
rect 4695 2806 4698 2814
rect 4702 2806 4703 2814
rect 4703 2806 4710 2814
rect 492 2796 500 2804
rect 908 2796 916 2804
rect 1228 2796 1236 2804
rect 1356 2796 1364 2804
rect 1196 2776 1204 2784
rect 1260 2776 1268 2784
rect 1484 2796 1492 2804
rect 1996 2796 2004 2804
rect 2156 2796 2164 2804
rect 3052 2796 3060 2804
rect 3788 2796 3796 2804
rect 3916 2796 3924 2804
rect 3948 2796 3956 2804
rect 4012 2796 4020 2804
rect 4076 2796 4084 2804
rect 4300 2796 4308 2804
rect 1516 2776 1524 2784
rect 1772 2776 1780 2784
rect 172 2756 180 2764
rect 940 2756 948 2764
rect 1228 2756 1236 2764
rect 1452 2756 1460 2764
rect 1708 2756 1716 2764
rect 2156 2756 2164 2764
rect 2348 2756 2356 2764
rect 2380 2756 2388 2764
rect 2732 2776 2740 2784
rect 3532 2776 3540 2784
rect 3756 2776 3764 2784
rect 4620 2776 4628 2784
rect 5324 2776 5332 2784
rect 5676 2776 5684 2784
rect 364 2736 372 2744
rect 556 2736 564 2744
rect 700 2716 708 2724
rect 1260 2736 1268 2744
rect 1100 2716 1108 2724
rect 1164 2716 1172 2724
rect 1388 2716 1396 2724
rect 1740 2736 1748 2744
rect 1964 2736 1972 2744
rect 1996 2736 2004 2744
rect 2732 2736 2740 2744
rect 3020 2760 3028 2768
rect 2764 2736 2772 2744
rect 3020 2732 3028 2740
rect 2124 2716 2132 2724
rect 2188 2716 2196 2724
rect 2860 2716 2868 2724
rect 3084 2716 3092 2724
rect 428 2696 436 2704
rect 620 2696 628 2704
rect 1004 2696 1012 2704
rect 364 2676 372 2684
rect 492 2676 500 2684
rect 524 2676 532 2684
rect 1676 2696 1684 2704
rect 1036 2676 1044 2684
rect 1068 2676 1076 2684
rect 1164 2676 1172 2684
rect 1260 2676 1268 2684
rect 1836 2696 1844 2704
rect 1996 2696 2004 2704
rect 2220 2696 2228 2704
rect 2700 2696 2708 2704
rect 2764 2696 2772 2704
rect 2988 2696 2996 2704
rect 3276 2736 3284 2744
rect 3308 2736 3316 2744
rect 3788 2736 3796 2744
rect 3820 2736 3828 2744
rect 4524 2756 4532 2764
rect 5932 2756 5940 2764
rect 3980 2736 3988 2744
rect 4492 2736 4500 2744
rect 5740 2736 5748 2744
rect 6156 2736 6164 2744
rect 3244 2716 3252 2724
rect 3404 2716 3412 2724
rect 3532 2716 3540 2724
rect 5580 2716 5588 2724
rect 5612 2716 5620 2724
rect 5708 2716 5716 2724
rect 3596 2696 3604 2704
rect 3628 2696 3636 2704
rect 1756 2676 1764 2684
rect 2188 2676 2196 2684
rect 2444 2676 2452 2684
rect 2476 2676 2484 2684
rect 460 2656 468 2664
rect 652 2656 660 2664
rect 716 2656 724 2664
rect 1164 2636 1172 2644
rect 1196 2656 1204 2664
rect 1420 2656 1428 2664
rect 1484 2636 1492 2644
rect 1772 2636 1780 2644
rect 1868 2656 1876 2664
rect 2252 2656 2260 2664
rect 1836 2636 1844 2644
rect 1964 2636 1972 2644
rect 2028 2636 2036 2644
rect 2348 2656 2356 2664
rect 2668 2656 2676 2664
rect 2732 2656 2740 2664
rect 2956 2676 2964 2684
rect 4108 2696 4116 2704
rect 4268 2696 4276 2704
rect 5708 2696 5716 2704
rect 6124 2716 6132 2724
rect 5900 2696 5908 2704
rect 6156 2696 6164 2704
rect 3276 2656 3284 2664
rect 3660 2656 3668 2664
rect 3724 2656 3732 2664
rect 3884 2656 3892 2664
rect 3948 2656 3956 2664
rect 3980 2656 3988 2664
rect 4172 2676 4180 2684
rect 4492 2676 4500 2684
rect 6188 2676 6196 2684
rect 5196 2656 5204 2664
rect 5484 2656 5492 2664
rect 5740 2656 5748 2664
rect 5932 2656 5940 2664
rect 6092 2656 6100 2664
rect 3308 2636 3316 2644
rect 5612 2636 5620 2644
rect 6124 2636 6132 2644
rect 6156 2636 6164 2644
rect 460 2616 468 2624
rect 684 2616 692 2624
rect 1068 2616 1076 2624
rect 1164 2616 1172 2624
rect 1868 2616 1876 2624
rect 2124 2616 2132 2624
rect 2252 2616 2260 2624
rect 2732 2616 2740 2624
rect 2764 2616 2772 2624
rect 716 2596 724 2604
rect 844 2596 852 2604
rect 1004 2596 1012 2604
rect 2220 2596 2228 2604
rect 2796 2596 2804 2604
rect 3468 2616 3476 2624
rect 3114 2606 3121 2614
rect 3121 2606 3122 2614
rect 3126 2606 3131 2614
rect 3131 2606 3133 2614
rect 3133 2606 3134 2614
rect 3138 2606 3141 2614
rect 3141 2606 3143 2614
rect 3143 2606 3146 2614
rect 3150 2606 3151 2614
rect 3151 2606 3158 2614
rect 2988 2596 2996 2604
rect 3436 2596 3444 2604
rect 3500 2596 3508 2604
rect 3628 2596 3636 2604
rect 3756 2616 3764 2624
rect 3916 2616 3924 2624
rect 4172 2616 4180 2624
rect 5324 2616 5332 2624
rect 5580 2616 5588 2624
rect 5804 2616 5812 2624
rect 108 2576 116 2584
rect 1484 2576 1492 2584
rect 1516 2576 1524 2584
rect 2476 2576 2484 2584
rect 3596 2576 3604 2584
rect 4044 2576 4052 2584
rect 4396 2596 4404 2604
rect 4492 2596 4500 2604
rect 4588 2596 4596 2604
rect 5932 2596 5940 2604
rect 6156 2596 6164 2604
rect 4620 2576 4628 2584
rect 4940 2576 4948 2584
rect 6028 2576 6036 2584
rect 204 2556 212 2564
rect 460 2556 468 2564
rect 716 2556 724 2564
rect 972 2556 980 2564
rect 1548 2556 1556 2564
rect 2524 2556 2532 2564
rect 140 2536 148 2544
rect 300 2536 308 2544
rect 524 2536 532 2544
rect 620 2536 628 2544
rect 652 2536 660 2544
rect 1292 2536 1300 2544
rect 1932 2536 1940 2544
rect 2028 2536 2036 2544
rect 2188 2536 2196 2544
rect 2316 2536 2324 2544
rect 2412 2536 2420 2544
rect 2636 2556 2644 2564
rect 2732 2556 2740 2564
rect 2956 2556 2964 2564
rect 3196 2556 3204 2564
rect 3404 2556 3412 2564
rect 3436 2556 3444 2564
rect 3820 2556 3828 2564
rect 3980 2556 3988 2564
rect 4108 2556 4116 2564
rect 5580 2556 5588 2564
rect 5772 2556 5780 2564
rect 2700 2536 2708 2544
rect 2892 2536 2900 2544
rect 3052 2536 3060 2544
rect 3084 2536 3092 2544
rect 3244 2536 3252 2544
rect 3532 2536 3540 2544
rect 3788 2536 3796 2544
rect 3916 2536 3924 2544
rect 4524 2536 4532 2544
rect 5260 2536 5268 2544
rect 5356 2536 5364 2544
rect 5644 2536 5652 2544
rect 12 2516 20 2524
rect 812 2516 820 2524
rect 1196 2516 1204 2524
rect 1356 2516 1364 2524
rect 2092 2516 2100 2524
rect 2524 2516 2532 2524
rect 3820 2516 3828 2524
rect 4076 2516 4084 2524
rect 4140 2516 4148 2524
rect 4172 2516 4180 2524
rect 5836 2516 5844 2524
rect 6060 2516 6068 2524
rect 6252 2536 6260 2544
rect 556 2496 564 2504
rect 1100 2496 1108 2504
rect 1324 2496 1332 2504
rect 1996 2496 2004 2504
rect 2060 2496 2068 2504
rect 492 2476 500 2484
rect 748 2476 756 2484
rect 1164 2476 1172 2484
rect 684 2456 692 2464
rect 716 2456 724 2464
rect 1420 2436 1428 2444
rect 1516 2476 1524 2484
rect 1676 2476 1684 2484
rect 1708 2476 1716 2484
rect 2156 2496 2164 2504
rect 2988 2496 2996 2504
rect 3084 2496 3092 2504
rect 3404 2496 3412 2504
rect 3436 2496 3444 2504
rect 2092 2476 2100 2484
rect 2396 2476 2404 2484
rect 2732 2476 2740 2484
rect 2924 2476 2932 2484
rect 3212 2476 3220 2484
rect 3980 2496 3988 2504
rect 4044 2496 4052 2504
rect 4268 2496 4276 2504
rect 4332 2496 4340 2504
rect 4428 2496 4436 2504
rect 5292 2496 5300 2504
rect 5804 2496 5812 2504
rect 5420 2476 5428 2484
rect 5772 2476 5780 2484
rect 3276 2456 3284 2464
rect 1452 2436 1460 2444
rect 2924 2436 2932 2444
rect 3020 2436 3028 2444
rect 3436 2456 3444 2464
rect 3692 2456 3700 2464
rect 3308 2436 3316 2444
rect 3884 2456 3892 2464
rect 4364 2456 4372 2464
rect 3948 2436 3956 2444
rect 4140 2436 4148 2444
rect 6028 2436 6036 2444
rect 684 2416 692 2424
rect 2060 2416 2068 2424
rect 3244 2416 3252 2424
rect 3756 2416 3764 2424
rect 5260 2416 5268 2424
rect 1578 2406 1585 2414
rect 1585 2406 1586 2414
rect 1590 2406 1595 2414
rect 1595 2406 1597 2414
rect 1597 2406 1598 2414
rect 1602 2406 1605 2414
rect 1605 2406 1607 2414
rect 1607 2406 1610 2414
rect 1614 2406 1615 2414
rect 1615 2406 1622 2414
rect 4666 2406 4673 2414
rect 4673 2406 4674 2414
rect 4678 2406 4683 2414
rect 4683 2406 4685 2414
rect 4685 2406 4686 2414
rect 4690 2406 4693 2414
rect 4693 2406 4695 2414
rect 4695 2406 4698 2414
rect 4702 2406 4703 2414
rect 4703 2406 4710 2414
rect 460 2396 468 2404
rect 1836 2396 1844 2404
rect 2092 2396 2100 2404
rect 2252 2396 2260 2404
rect 2284 2396 2292 2404
rect 2316 2396 2324 2404
rect 2636 2396 2644 2404
rect 3196 2396 3204 2404
rect 76 2376 84 2384
rect 844 2376 852 2384
rect 780 2356 788 2364
rect 1516 2356 1524 2364
rect 1644 2356 1652 2364
rect 2380 2376 2388 2384
rect 2860 2376 2868 2384
rect 2988 2376 2996 2384
rect 3052 2376 3060 2384
rect 3468 2396 3476 2404
rect 4044 2396 4052 2404
rect 5804 2396 5812 2404
rect 3308 2376 3316 2384
rect 4268 2376 4276 2384
rect 2060 2356 2068 2364
rect 2220 2356 2228 2364
rect 6252 2356 6260 2364
rect 428 2336 436 2344
rect 684 2336 692 2344
rect 1004 2336 1012 2344
rect 1292 2336 1300 2344
rect 1388 2336 1396 2344
rect 1452 2336 1460 2344
rect 2124 2336 2132 2344
rect 2892 2336 2900 2344
rect 780 2316 788 2324
rect 1644 2316 1652 2324
rect 2220 2316 2228 2324
rect 2524 2316 2532 2324
rect 2988 2316 2996 2324
rect 3884 2336 3892 2344
rect 4332 2336 4340 2344
rect 4588 2336 4596 2344
rect 5324 2336 5332 2344
rect 5676 2336 5684 2344
rect 5772 2336 5780 2344
rect 6060 2336 6068 2344
rect 12 2296 20 2304
rect 524 2296 532 2304
rect 2252 2296 2260 2304
rect 428 2256 436 2264
rect 972 2276 980 2284
rect 1356 2276 1364 2284
rect 1740 2276 1748 2284
rect 1964 2276 1972 2284
rect 2092 2256 2100 2264
rect 2188 2256 2196 2264
rect 2380 2296 2388 2304
rect 2476 2296 2484 2304
rect 2540 2296 2548 2304
rect 2572 2276 2580 2284
rect 2604 2280 2612 2288
rect 2636 2276 2644 2284
rect 2764 2296 2772 2304
rect 3020 2296 3028 2304
rect 3532 2296 3540 2304
rect 3628 2296 3636 2304
rect 3788 2296 3796 2304
rect 4204 2296 4212 2304
rect 4492 2296 4500 2304
rect 5068 2296 5076 2304
rect 5676 2296 5684 2304
rect 2860 2276 2868 2284
rect 2892 2276 2900 2284
rect 3052 2276 3060 2284
rect 3244 2276 3252 2284
rect 3372 2276 3380 2284
rect 2316 2256 2324 2264
rect 2508 2256 2516 2264
rect 2604 2252 2612 2260
rect 2764 2256 2772 2264
rect 2924 2256 2932 2264
rect 2956 2256 2964 2264
rect 780 2236 788 2244
rect 1868 2236 1876 2244
rect 3180 2256 3188 2264
rect 3276 2256 3284 2264
rect 3436 2256 3444 2264
rect 3596 2276 3604 2284
rect 3692 2276 3700 2284
rect 3756 2276 3764 2284
rect 396 2216 404 2224
rect 844 2216 852 2224
rect 1804 2216 1812 2224
rect 3788 2256 3796 2264
rect 4140 2276 4148 2284
rect 5836 2276 5844 2284
rect 5932 2276 5940 2284
rect 3916 2256 3924 2264
rect 4236 2256 4244 2264
rect 5804 2256 5812 2264
rect 3628 2236 3636 2244
rect 4108 2236 4116 2244
rect 4460 2236 4468 2244
rect 3308 2216 3316 2224
rect 5676 2216 5684 2224
rect 3114 2206 3121 2214
rect 3121 2206 3122 2214
rect 3126 2206 3131 2214
rect 3131 2206 3133 2214
rect 3133 2206 3134 2214
rect 3138 2206 3141 2214
rect 3141 2206 3143 2214
rect 3143 2206 3146 2214
rect 3150 2206 3151 2214
rect 3151 2206 3158 2214
rect 428 2196 436 2204
rect 652 2196 660 2204
rect 748 2196 756 2204
rect 1068 2196 1076 2204
rect 1868 2196 1876 2204
rect 2028 2196 2036 2204
rect 2348 2196 2356 2204
rect 492 2176 500 2184
rect 1420 2176 1428 2184
rect 1740 2176 1748 2184
rect 1836 2176 1844 2184
rect 1932 2176 1940 2184
rect 652 2156 660 2164
rect 844 2156 852 2164
rect 1004 2156 1012 2164
rect 588 2136 596 2144
rect 172 2116 180 2124
rect 396 2116 404 2124
rect 620 2116 628 2124
rect 652 2116 660 2124
rect 1036 2136 1044 2144
rect 1260 2136 1268 2144
rect 1388 2136 1396 2144
rect 1708 2156 1716 2164
rect 1772 2156 1780 2164
rect 1868 2156 1876 2164
rect 2252 2176 2260 2184
rect 2284 2176 2292 2184
rect 2396 2196 2404 2204
rect 2476 2196 2484 2204
rect 2668 2196 2676 2204
rect 3052 2196 3060 2204
rect 3468 2196 3476 2204
rect 3980 2196 3988 2204
rect 4300 2196 4308 2204
rect 4364 2196 4372 2204
rect 5036 2196 5044 2204
rect 2124 2156 2132 2164
rect 1644 2136 1652 2144
rect 1196 2116 1204 2124
rect 1676 2136 1684 2144
rect 1932 2136 1940 2144
rect 2348 2156 2356 2164
rect 2540 2156 2548 2164
rect 2636 2156 2644 2164
rect 2668 2156 2676 2164
rect 3404 2176 3412 2184
rect 3308 2156 3316 2164
rect 3532 2156 3540 2164
rect 3916 2176 3924 2184
rect 4172 2176 4180 2184
rect 4236 2176 4244 2184
rect 4876 2176 4884 2184
rect 5132 2176 5140 2184
rect 5804 2176 5812 2184
rect 5836 2176 5844 2184
rect 2156 2136 2164 2144
rect 2572 2136 2580 2144
rect 2988 2136 2996 2144
rect 1708 2116 1716 2124
rect 1740 2116 1748 2124
rect 1804 2116 1812 2124
rect 364 2096 372 2104
rect 556 2076 564 2084
rect 588 2076 596 2084
rect 1228 2096 1236 2104
rect 3852 2136 3860 2144
rect 4268 2156 4276 2164
rect 4588 2156 4596 2164
rect 4332 2136 4340 2144
rect 4396 2136 4404 2144
rect 1996 2096 2004 2104
rect 2060 2096 2068 2104
rect 2156 2096 2164 2104
rect 2220 2096 2228 2104
rect 2476 2096 2484 2104
rect 2508 2096 2516 2104
rect 2732 2096 2740 2104
rect 3244 2096 3252 2104
rect 3404 2096 3412 2104
rect 6028 2136 6036 2144
rect 4620 2116 4628 2124
rect 4844 2116 4852 2124
rect 4940 2116 4948 2124
rect 5036 2116 5044 2124
rect 3852 2096 3860 2104
rect 4108 2096 4116 2104
rect 4300 2096 4308 2104
rect 5004 2096 5012 2104
rect 5132 2096 5140 2104
rect 1068 2076 1076 2084
rect 1100 2076 1108 2084
rect 1388 2076 1396 2084
rect 1804 2076 1812 2084
rect 1980 2076 1988 2084
rect 2860 2076 2868 2084
rect 2988 2076 2996 2084
rect 3180 2076 3188 2084
rect 3500 2076 3508 2084
rect 3660 2076 3668 2084
rect 4588 2076 4596 2084
rect 4620 2076 4628 2084
rect 6028 2076 6036 2084
rect 1324 2056 1332 2064
rect 1644 2056 1652 2064
rect 1772 2056 1780 2064
rect 2956 2056 2964 2064
rect 3020 2056 3028 2064
rect 3340 2056 3348 2064
rect 3916 2056 3924 2064
rect 3948 2056 3956 2064
rect 4460 2056 4468 2064
rect 6092 2056 6100 2064
rect 2540 2036 2548 2044
rect 4044 2036 4052 2044
rect 4172 2036 4180 2044
rect 4236 2036 4244 2044
rect 4364 2036 4372 2044
rect 4780 2036 4788 2044
rect 4844 2036 4852 2044
rect 5612 2036 5620 2044
rect 492 2016 500 2024
rect 908 2016 916 2024
rect 940 2016 948 2024
rect 1068 2016 1076 2024
rect 1388 2016 1396 2024
rect 2476 2016 2484 2024
rect 2604 2016 2612 2024
rect 2636 2016 2644 2024
rect 2764 2016 2772 2024
rect 2796 2016 2804 2024
rect 1578 2006 1585 2014
rect 1585 2006 1586 2014
rect 1590 2006 1595 2014
rect 1595 2006 1597 2014
rect 1597 2006 1598 2014
rect 1602 2006 1605 2014
rect 1605 2006 1607 2014
rect 1607 2006 1610 2014
rect 1614 2006 1615 2014
rect 1615 2006 1622 2014
rect 1132 1996 1140 2004
rect 1196 1996 1204 2004
rect 1356 1996 1364 2004
rect 1404 1996 1412 2004
rect 1676 1996 1684 2004
rect 1708 1996 1716 2004
rect 1964 1996 1972 2004
rect 2508 1996 2516 2004
rect 2892 1996 2900 2004
rect 3212 1996 3220 2004
rect 3660 2016 3668 2024
rect 4666 2006 4673 2014
rect 4673 2006 4674 2014
rect 4678 2006 4683 2014
rect 4683 2006 4685 2014
rect 4685 2006 4686 2014
rect 4690 2006 4693 2014
rect 4693 2006 4695 2014
rect 4695 2006 4698 2014
rect 4702 2006 4703 2014
rect 4703 2006 4710 2014
rect 1036 1976 1044 1984
rect 1868 1976 1876 1984
rect 1996 1976 2004 1984
rect 2092 1976 2100 1984
rect 2252 1976 2260 1984
rect 396 1956 404 1964
rect 492 1956 500 1964
rect 556 1936 564 1944
rect 652 1936 660 1944
rect 1388 1956 1396 1964
rect 1420 1956 1428 1964
rect 1484 1936 1492 1944
rect 3340 1996 3348 2004
rect 3372 1996 3380 2004
rect 3404 1996 3412 2004
rect 3532 1996 3540 2004
rect 3596 1996 3604 2004
rect 3756 1976 3764 1984
rect 3980 1996 3988 2004
rect 4140 1996 4148 2004
rect 3948 1976 3956 1984
rect 5004 1996 5012 2004
rect 6092 1996 6100 2004
rect 5420 1976 5428 1984
rect 2924 1956 2932 1964
rect 3020 1956 3028 1964
rect 3276 1956 3284 1964
rect 3308 1956 3316 1964
rect 4396 1956 4404 1964
rect 4588 1956 4596 1964
rect 1900 1936 1908 1944
rect 1932 1936 1940 1944
rect 620 1916 628 1924
rect 1292 1916 1300 1924
rect 1324 1916 1332 1924
rect 108 1896 116 1904
rect 364 1896 372 1904
rect 1740 1916 1748 1924
rect 2124 1936 2132 1944
rect 2220 1936 2228 1944
rect 3212 1936 3220 1944
rect 3660 1936 3668 1944
rect 5356 1936 5364 1944
rect 5740 1936 5748 1944
rect 2156 1916 2164 1924
rect 2412 1916 2420 1924
rect 2924 1920 2932 1928
rect 2956 1916 2964 1924
rect 3308 1916 3316 1924
rect 3356 1916 3364 1924
rect 1868 1896 1876 1904
rect 1932 1896 1940 1904
rect 2028 1896 2036 1904
rect 2060 1896 2068 1904
rect 2188 1896 2196 1904
rect 2828 1896 2836 1904
rect 2924 1896 2932 1900
rect 3468 1916 3476 1924
rect 3820 1916 3828 1924
rect 3852 1916 3860 1924
rect 4140 1916 4148 1924
rect 3532 1896 3540 1904
rect 2924 1892 2932 1896
rect 1132 1876 1140 1884
rect 1292 1876 1300 1884
rect 1484 1876 1492 1884
rect 172 1856 180 1864
rect 876 1856 884 1864
rect 1228 1856 1236 1864
rect 844 1836 852 1844
rect 1708 1876 1716 1884
rect 2092 1876 2100 1884
rect 2156 1876 2164 1884
rect 2332 1876 2340 1884
rect 1420 1836 1428 1844
rect 1068 1816 1076 1824
rect 1164 1816 1172 1824
rect 1292 1816 1300 1824
rect 1324 1816 1332 1824
rect 1356 1816 1364 1824
rect 1388 1816 1396 1824
rect 1676 1856 1684 1864
rect 1836 1856 1844 1864
rect 1548 1816 1556 1824
rect 1644 1816 1652 1824
rect 1900 1856 1908 1864
rect 1996 1856 2004 1864
rect 2252 1856 2260 1864
rect 2380 1856 2388 1864
rect 2716 1876 2724 1884
rect 2764 1876 2772 1884
rect 2892 1876 2900 1884
rect 3052 1876 3060 1884
rect 3404 1876 3412 1884
rect 3564 1876 3572 1884
rect 3884 1876 3892 1884
rect 3980 1876 3988 1884
rect 4044 1896 4052 1904
rect 4844 1916 4852 1924
rect 4908 1916 4916 1924
rect 5068 1916 5076 1924
rect 5100 1916 5108 1924
rect 5548 1916 5556 1924
rect 4204 1896 4212 1904
rect 4524 1896 4532 1904
rect 4620 1896 4628 1904
rect 4876 1896 4884 1904
rect 5292 1896 5300 1904
rect 5708 1896 5716 1904
rect 5324 1876 5332 1884
rect 5452 1876 5460 1884
rect 6252 1876 6260 1884
rect 1740 1816 1748 1824
rect 1836 1816 1844 1824
rect 2092 1836 2100 1844
rect 2284 1836 2292 1844
rect 2156 1816 2164 1824
rect 2604 1836 2612 1844
rect 2700 1856 2708 1864
rect 3180 1856 3188 1864
rect 2316 1816 2324 1824
rect 2380 1816 2388 1824
rect 2444 1816 2452 1824
rect 2572 1816 2580 1824
rect 2668 1816 2676 1824
rect 2732 1836 2740 1844
rect 3020 1836 3028 1844
rect 3308 1856 3316 1864
rect 3340 1856 3348 1864
rect 4140 1856 4148 1864
rect 3372 1836 3380 1844
rect 3244 1816 3252 1824
rect 3276 1816 3284 1824
rect 3628 1836 3636 1844
rect 3692 1836 3700 1844
rect 4620 1836 4628 1844
rect 4780 1836 4788 1844
rect 4844 1856 4852 1864
rect 5100 1856 5108 1864
rect 5708 1856 5716 1864
rect 5932 1856 5940 1864
rect 3852 1816 3860 1824
rect 2124 1796 2132 1804
rect 2188 1796 2196 1804
rect 2348 1796 2356 1804
rect 2540 1796 2548 1804
rect 2956 1800 2964 1808
rect 3114 1806 3121 1814
rect 3121 1806 3122 1814
rect 3126 1806 3131 1814
rect 3131 1806 3133 1814
rect 3133 1806 3134 1814
rect 3138 1806 3141 1814
rect 3141 1806 3143 1814
rect 3143 1806 3146 1814
rect 3150 1806 3151 1814
rect 3151 1806 3158 1814
rect 3020 1796 3028 1804
rect 3212 1796 3220 1804
rect 3532 1796 3540 1804
rect 3692 1796 3700 1804
rect 3724 1796 3732 1804
rect 4844 1816 4852 1824
rect 4908 1816 4916 1824
rect 6028 1816 6036 1824
rect 4204 1796 4212 1804
rect 4332 1796 4340 1804
rect 2252 1776 2260 1784
rect 2284 1776 2292 1784
rect 2476 1780 2484 1788
rect 2700 1776 2708 1784
rect 2956 1772 2964 1780
rect 4876 1776 4884 1784
rect 5004 1776 5012 1784
rect 5516 1776 5524 1784
rect 76 1756 84 1764
rect 1100 1756 1108 1764
rect 1516 1756 1524 1764
rect 812 1736 820 1744
rect 1996 1756 2004 1764
rect 2060 1736 2068 1744
rect 2156 1736 2164 1744
rect 2316 1736 2324 1744
rect 620 1716 628 1724
rect 1324 1716 1332 1724
rect 1420 1716 1428 1724
rect 1708 1716 1716 1724
rect 1836 1716 1844 1724
rect 1900 1716 1908 1724
rect 1964 1716 1972 1724
rect 2284 1716 2292 1724
rect 2348 1736 2356 1744
rect 2476 1752 2484 1760
rect 3084 1756 3092 1764
rect 3212 1756 3220 1764
rect 3724 1756 3732 1764
rect 3788 1756 3796 1764
rect 3996 1756 4004 1764
rect 2700 1736 2708 1744
rect 2796 1736 2804 1744
rect 2956 1736 2964 1744
rect 2988 1736 2996 1744
rect 3500 1736 3508 1744
rect 4268 1736 4276 1744
rect 4332 1736 4340 1744
rect 4428 1736 4436 1744
rect 4556 1736 4564 1744
rect 4972 1736 4980 1744
rect 5324 1736 5332 1744
rect 5836 1736 5844 1744
rect 2444 1716 2452 1724
rect 3372 1716 3380 1724
rect 3468 1716 3476 1724
rect 3756 1716 3764 1724
rect 4268 1716 4276 1724
rect 5612 1716 5620 1724
rect 6028 1716 6036 1724
rect 588 1696 596 1704
rect 1036 1696 1044 1704
rect 1068 1696 1076 1704
rect 1196 1696 1204 1704
rect 460 1676 468 1684
rect 1868 1696 1876 1704
rect 2156 1696 2164 1704
rect 2700 1696 2708 1704
rect 2892 1696 2900 1704
rect 3820 1696 3828 1704
rect 1548 1676 1556 1684
rect 1996 1676 2004 1684
rect 2220 1676 2228 1684
rect 2380 1676 2388 1684
rect 2540 1676 2548 1684
rect 908 1656 916 1664
rect 1004 1636 1012 1644
rect 1132 1656 1140 1664
rect 1260 1656 1268 1664
rect 1388 1656 1396 1664
rect 2060 1656 2068 1664
rect 2636 1676 2644 1684
rect 2764 1676 2772 1684
rect 2828 1676 2836 1684
rect 2924 1676 2932 1684
rect 3244 1676 3252 1684
rect 4108 1696 4116 1704
rect 4172 1696 4180 1704
rect 4300 1696 4308 1704
rect 4428 1696 4436 1704
rect 4492 1696 4500 1704
rect 5452 1696 5460 1704
rect 6252 1696 6260 1704
rect 2700 1656 2708 1664
rect 5708 1676 5716 1684
rect 4748 1656 4756 1664
rect 4876 1656 4884 1664
rect 5452 1656 5460 1664
rect 5612 1656 5620 1664
rect 1068 1636 1076 1644
rect 1996 1636 2004 1644
rect 2540 1636 2548 1644
rect 3404 1636 3412 1644
rect 5036 1636 5044 1644
rect 5484 1636 5492 1644
rect 1100 1616 1108 1624
rect 1260 1616 1268 1624
rect 1356 1616 1364 1624
rect 2796 1616 2804 1624
rect 2892 1616 2900 1624
rect 4044 1616 4052 1624
rect 4268 1616 4276 1624
rect 1578 1606 1585 1614
rect 1585 1606 1586 1614
rect 1590 1606 1595 1614
rect 1595 1606 1597 1614
rect 1597 1606 1598 1614
rect 1602 1606 1605 1614
rect 1605 1606 1607 1614
rect 1607 1606 1610 1614
rect 1614 1606 1615 1614
rect 1615 1606 1622 1614
rect 5388 1616 5396 1624
rect 4666 1606 4673 1614
rect 4673 1606 4674 1614
rect 4678 1606 4683 1614
rect 4683 1606 4685 1614
rect 4685 1606 4686 1614
rect 4690 1606 4693 1614
rect 4693 1606 4695 1614
rect 4695 1606 4698 1614
rect 4702 1606 4703 1614
rect 4703 1606 4710 1614
rect 972 1596 980 1604
rect 1004 1576 1012 1584
rect 1356 1576 1364 1584
rect 1916 1596 1924 1604
rect 2572 1596 2580 1604
rect 3532 1596 3540 1604
rect 3756 1596 3764 1604
rect 3916 1596 3924 1604
rect 4236 1596 4244 1604
rect 4300 1596 4308 1604
rect 4588 1596 4596 1604
rect 1868 1576 1876 1584
rect 1964 1576 1972 1584
rect 3468 1576 3476 1584
rect 4012 1576 4020 1584
rect 4332 1576 4340 1584
rect 4492 1576 4500 1584
rect 5484 1576 5492 1584
rect 492 1556 500 1564
rect 876 1556 884 1564
rect 940 1536 948 1544
rect 1100 1536 1108 1544
rect 1548 1536 1556 1544
rect 1644 1536 1652 1544
rect 428 1516 436 1524
rect 236 1496 244 1504
rect 524 1496 532 1504
rect 556 1496 564 1504
rect 716 1496 724 1504
rect 364 1476 372 1484
rect 812 1516 820 1524
rect 780 1496 788 1504
rect 1132 1516 1140 1524
rect 1228 1516 1236 1524
rect 1292 1516 1300 1524
rect 1484 1516 1492 1524
rect 1740 1536 1748 1544
rect 1836 1536 1844 1544
rect 2124 1536 2132 1544
rect 2284 1536 2292 1544
rect 2380 1536 2388 1544
rect 3660 1556 3668 1564
rect 3788 1556 3796 1564
rect 3916 1556 3924 1564
rect 4204 1556 4212 1564
rect 4556 1556 4564 1564
rect 4588 1556 4596 1564
rect 2732 1536 2740 1544
rect 2764 1536 2772 1544
rect 3564 1536 3572 1544
rect 4396 1536 4404 1544
rect 4460 1536 4468 1544
rect 1932 1516 1940 1524
rect 2092 1516 2100 1524
rect 2316 1516 2324 1524
rect 2412 1516 2420 1524
rect 3020 1516 3028 1524
rect 3084 1516 3092 1524
rect 3308 1516 3316 1524
rect 1260 1476 1268 1484
rect 1452 1496 1460 1504
rect 1644 1496 1652 1504
rect 2060 1496 2068 1504
rect 2796 1496 2804 1504
rect 812 1456 820 1464
rect 1004 1456 1012 1464
rect 1196 1456 1204 1464
rect 1420 1456 1428 1464
rect 1868 1476 1876 1484
rect 2092 1476 2100 1484
rect 2252 1476 2260 1484
rect 2284 1476 2292 1484
rect 2476 1476 2484 1484
rect 2156 1456 2164 1464
rect 2188 1456 2196 1464
rect 2508 1456 2516 1464
rect 2572 1456 2580 1464
rect 2700 1476 2708 1484
rect 2924 1476 2932 1484
rect 3372 1496 3380 1504
rect 4300 1496 4308 1504
rect 5164 1556 5172 1564
rect 5772 1556 5780 1564
rect 5196 1536 5204 1544
rect 5260 1536 5268 1544
rect 5772 1516 5780 1524
rect 6252 1536 6260 1544
rect 4460 1500 4468 1508
rect 4812 1496 4820 1504
rect 4940 1496 4948 1504
rect 5516 1496 5524 1504
rect 5580 1496 5588 1504
rect 5708 1496 5716 1504
rect 6060 1496 6068 1504
rect 3212 1476 3220 1484
rect 3404 1476 3412 1484
rect 3468 1476 3476 1484
rect 4044 1476 4052 1484
rect 4268 1476 4276 1484
rect 4460 1472 4468 1480
rect 4524 1476 4532 1484
rect 2764 1456 2772 1464
rect 2796 1456 2804 1464
rect 3372 1456 3380 1464
rect 3532 1456 3540 1464
rect 4588 1456 4596 1464
rect 4748 1476 4756 1484
rect 5260 1476 5268 1484
rect 5324 1476 5332 1484
rect 5996 1476 6004 1484
rect 6252 1496 6260 1504
rect 748 1416 756 1424
rect 1228 1436 1236 1444
rect 1260 1436 1268 1444
rect 1772 1436 1780 1444
rect 2060 1436 2068 1444
rect 844 1416 852 1424
rect 1004 1416 1012 1424
rect 1164 1416 1172 1424
rect 1356 1416 1364 1424
rect 1516 1416 1524 1424
rect 3020 1436 3028 1444
rect 3308 1436 3316 1444
rect 3436 1436 3444 1444
rect 3788 1436 3796 1444
rect 4204 1436 4212 1444
rect 4556 1436 4564 1444
rect 5132 1456 5140 1464
rect 5580 1456 5588 1464
rect 5836 1456 5844 1464
rect 4876 1436 4884 1444
rect 5484 1436 5492 1444
rect 5932 1436 5940 1444
rect 2252 1416 2260 1424
rect 2444 1416 2452 1424
rect 2508 1416 2516 1424
rect 3212 1416 3220 1424
rect 3404 1416 3412 1424
rect 3660 1416 3668 1424
rect 4140 1416 4148 1424
rect 6028 1416 6036 1424
rect 3114 1406 3121 1414
rect 3121 1406 3122 1414
rect 3126 1406 3131 1414
rect 3131 1406 3133 1414
rect 3133 1406 3134 1414
rect 3138 1406 3141 1414
rect 3141 1406 3143 1414
rect 3143 1406 3146 1414
rect 3150 1406 3151 1414
rect 3151 1406 3158 1414
rect 908 1396 916 1404
rect 1100 1396 1108 1404
rect 1676 1396 1684 1404
rect 1836 1396 1844 1404
rect 844 1376 852 1384
rect 1228 1376 1236 1384
rect 2828 1396 2836 1404
rect 4076 1396 4084 1404
rect 4236 1396 4244 1404
rect 4268 1396 4276 1404
rect 4620 1396 4628 1404
rect 4844 1396 4852 1404
rect 5772 1396 5780 1404
rect 5932 1396 5940 1404
rect 5964 1396 5972 1404
rect 268 1336 276 1344
rect 300 1336 308 1344
rect 876 1336 884 1344
rect 940 1356 948 1364
rect 1356 1356 1364 1364
rect 1388 1356 1396 1364
rect 1420 1356 1428 1364
rect 1484 1356 1492 1364
rect 1548 1356 1556 1364
rect 1836 1356 1844 1364
rect 2188 1356 2196 1364
rect 2252 1356 2260 1364
rect 2316 1356 2324 1364
rect 3020 1376 3028 1384
rect 3212 1376 3220 1384
rect 3532 1376 3540 1384
rect 3980 1376 3988 1384
rect 4108 1376 4116 1384
rect 4332 1376 4340 1384
rect 4492 1376 4500 1384
rect 172 1316 180 1324
rect 716 1316 724 1324
rect 1164 1316 1172 1324
rect 1292 1316 1300 1324
rect 1484 1316 1492 1324
rect 1740 1316 1748 1324
rect 1964 1316 1972 1324
rect 2092 1316 2100 1324
rect 2348 1336 2356 1344
rect 2444 1316 2452 1324
rect 2572 1316 2580 1324
rect 2700 1316 2708 1324
rect 2764 1316 2772 1324
rect 3020 1336 3028 1344
rect 3372 1336 3380 1344
rect 3436 1336 3444 1344
rect 3628 1356 3636 1364
rect 3660 1356 3668 1364
rect 4076 1356 4084 1364
rect 5836 1356 5844 1364
rect 6028 1356 6036 1364
rect 3788 1336 3796 1344
rect 3884 1336 3892 1344
rect 4108 1336 4116 1344
rect 4140 1336 4148 1344
rect 5036 1336 5044 1344
rect 5964 1336 5972 1344
rect 5996 1336 6004 1344
rect 2844 1316 2852 1324
rect 2988 1316 2996 1324
rect 3180 1316 3188 1324
rect 3500 1316 3508 1324
rect 5228 1316 5236 1324
rect 5356 1316 5364 1324
rect 5516 1316 5524 1324
rect 1004 1296 1012 1304
rect 1068 1296 1076 1304
rect 1356 1296 1364 1304
rect 1708 1296 1716 1304
rect 1164 1276 1172 1284
rect 1260 1276 1268 1284
rect 2028 1296 2036 1304
rect 2060 1296 2068 1304
rect 2412 1296 2420 1304
rect 3052 1296 3060 1304
rect 3276 1296 3284 1304
rect 3372 1296 3380 1304
rect 3468 1296 3476 1304
rect 3916 1296 3924 1304
rect 4524 1296 4532 1304
rect 5004 1296 5012 1304
rect 1036 1256 1044 1264
rect 1484 1256 1492 1264
rect 1964 1276 1972 1284
rect 2124 1276 2132 1284
rect 2348 1276 2356 1284
rect 2380 1276 2388 1284
rect 2636 1276 2644 1284
rect 2796 1276 2804 1284
rect 2828 1276 2836 1284
rect 2892 1276 2900 1284
rect 3500 1276 3508 1284
rect 3660 1276 3668 1284
rect 3852 1276 3860 1284
rect 4556 1276 4564 1284
rect 4588 1276 4596 1284
rect 4780 1276 4788 1284
rect 4876 1276 4884 1284
rect 4908 1276 4916 1284
rect 5292 1276 5300 1284
rect 5452 1276 5460 1284
rect 5612 1316 5620 1324
rect 2092 1256 2100 1264
rect 3244 1256 3252 1264
rect 3276 1256 3284 1264
rect 3404 1256 3412 1264
rect 3596 1256 3604 1264
rect 4332 1256 4340 1264
rect 5036 1256 5044 1264
rect 1516 1216 1524 1224
rect 1676 1216 1684 1224
rect 2284 1236 2292 1244
rect 2348 1236 2356 1244
rect 2604 1236 2612 1244
rect 5100 1236 5108 1244
rect 5292 1236 5300 1244
rect 6060 1276 6068 1284
rect 972 1196 980 1204
rect 1004 1196 1012 1204
rect 1292 1196 1300 1204
rect 1578 1206 1585 1214
rect 1585 1206 1586 1214
rect 1590 1206 1595 1214
rect 1595 1206 1597 1214
rect 1597 1206 1598 1214
rect 1602 1206 1605 1214
rect 1605 1206 1607 1214
rect 1607 1206 1610 1214
rect 1614 1206 1615 1214
rect 1615 1206 1622 1214
rect 76 1176 84 1184
rect 940 1176 948 1184
rect 1068 1176 1076 1184
rect 1132 1176 1140 1184
rect 1164 1176 1172 1184
rect 1804 1196 1812 1204
rect 2220 1196 2228 1204
rect 2252 1196 2260 1204
rect 2284 1196 2292 1204
rect 2316 1216 2324 1224
rect 4460 1216 4468 1224
rect 4492 1216 4500 1224
rect 4588 1216 4596 1224
rect 5164 1216 5172 1224
rect 5484 1216 5492 1224
rect 5612 1216 5620 1224
rect 6060 1216 6068 1224
rect 4666 1206 4673 1214
rect 4673 1206 4674 1214
rect 4678 1206 4683 1214
rect 4683 1206 4685 1214
rect 4685 1206 4686 1214
rect 4690 1206 4693 1214
rect 4693 1206 4695 1214
rect 4695 1206 4698 1214
rect 4702 1206 4703 1214
rect 4703 1206 4710 1214
rect 2732 1196 2740 1204
rect 2156 1176 2164 1184
rect 2316 1176 2324 1184
rect 2700 1176 2708 1184
rect 3724 1196 3732 1204
rect 4556 1196 4564 1204
rect 4748 1196 4756 1204
rect 2796 1176 2804 1184
rect 3212 1176 3220 1184
rect 3756 1176 3764 1184
rect 5772 1196 5780 1204
rect 6220 1196 6228 1204
rect 748 1156 756 1164
rect 2636 1156 2644 1164
rect 3052 1156 3060 1164
rect 4108 1156 4116 1164
rect 4300 1156 4308 1164
rect 4428 1156 4436 1164
rect 5260 1156 5268 1164
rect 5836 1156 5844 1164
rect 6220 1156 6228 1164
rect 716 1136 724 1144
rect 812 1136 820 1144
rect 844 1136 852 1144
rect 1676 1136 1684 1144
rect 172 1116 180 1124
rect 940 1116 948 1124
rect 972 1116 980 1124
rect 1452 1116 1460 1124
rect 12 1096 20 1104
rect 268 1096 276 1104
rect 908 1096 916 1104
rect 1260 1096 1268 1104
rect 1708 1116 1716 1124
rect 1836 1116 1844 1124
rect 3372 1136 3380 1144
rect 4076 1136 4084 1144
rect 4556 1136 4564 1144
rect 524 1076 532 1084
rect 300 1056 308 1064
rect 652 1056 660 1064
rect 780 1056 788 1064
rect 1100 1076 1108 1084
rect 1484 1076 1492 1084
rect 2220 1116 2228 1124
rect 2540 1116 2548 1124
rect 2604 1116 2612 1124
rect 3180 1116 3188 1124
rect 3532 1116 3540 1124
rect 4428 1116 4436 1124
rect 4460 1116 4468 1124
rect 4524 1116 4532 1124
rect 1964 1096 1972 1104
rect 2668 1096 2676 1104
rect 3340 1096 3348 1104
rect 3564 1096 3572 1104
rect 4172 1096 4180 1104
rect 4556 1096 4564 1104
rect 4620 1116 4628 1124
rect 4748 1116 4756 1124
rect 4844 1116 4852 1124
rect 5132 1116 5140 1124
rect 5964 1136 5972 1144
rect 5836 1116 5844 1124
rect 1804 1076 1812 1084
rect 1868 1076 1876 1084
rect 1932 1076 1940 1084
rect 2188 1076 2196 1084
rect 2220 1076 2228 1084
rect 1356 1036 1364 1044
rect 2540 1076 2548 1084
rect 2924 1076 2932 1084
rect 3084 1076 3092 1084
rect 3532 1076 3540 1084
rect 3820 1076 3828 1084
rect 4364 1076 4372 1084
rect 4588 1076 4596 1084
rect 4972 1096 4980 1104
rect 5548 1096 5556 1104
rect 6188 1116 6196 1124
rect 5868 1096 5876 1104
rect 4780 1076 4788 1084
rect 5068 1076 5076 1084
rect 5324 1076 5332 1084
rect 5516 1076 5524 1084
rect 5964 1076 5972 1084
rect 5996 1076 6004 1084
rect 2636 1056 2644 1064
rect 2892 1056 2900 1064
rect 3244 1056 3252 1064
rect 4204 1056 4212 1064
rect 4844 1056 4852 1064
rect 4876 1056 4884 1064
rect 5420 1056 5428 1064
rect 5484 1056 5492 1064
rect 1644 1036 1652 1044
rect 1708 1036 1716 1044
rect 76 1016 84 1024
rect 428 996 436 1004
rect 716 996 724 1004
rect 812 996 820 1004
rect 844 996 852 1004
rect 876 996 884 1004
rect 988 996 996 1004
rect 1068 996 1076 1004
rect 1836 1036 1844 1044
rect 1964 1036 1972 1044
rect 2604 1036 2612 1044
rect 3916 1036 3924 1044
rect 4332 1036 4340 1044
rect 4460 1036 4468 1044
rect 5228 1036 5236 1044
rect 2316 1016 2324 1024
rect 2348 1016 2356 1024
rect 2380 1016 2388 1024
rect 3114 1006 3121 1014
rect 3121 1006 3122 1014
rect 3126 1006 3131 1014
rect 3131 1006 3133 1014
rect 3133 1006 3134 1014
rect 3138 1006 3141 1014
rect 3141 1006 3143 1014
rect 3143 1006 3146 1014
rect 3150 1006 3151 1014
rect 3151 1006 3158 1014
rect 1164 996 1172 1004
rect 1196 996 1204 1004
rect 1516 996 1524 1004
rect 1548 996 1556 1004
rect 1964 996 1972 1004
rect 2220 996 2228 1004
rect 2412 996 2420 1004
rect 2540 996 2548 1004
rect 268 976 276 984
rect 1132 976 1140 984
rect 1452 976 1460 984
rect 2092 976 2100 984
rect 2124 976 2132 984
rect 2316 976 2324 984
rect 2764 976 2772 984
rect 2860 976 2868 984
rect 3244 976 3252 984
rect 3340 976 3348 984
rect 3500 996 3508 1004
rect 4268 1016 4276 1024
rect 4364 1016 4372 1024
rect 4556 1016 4564 1024
rect 5068 1016 5076 1024
rect 5388 1016 5396 1024
rect 5612 1016 5620 1024
rect 5836 1016 5844 1024
rect 5868 1016 5876 1024
rect 4204 996 4212 1004
rect 4332 996 4340 1004
rect 4780 996 4788 1004
rect 4844 996 4852 1004
rect 5036 996 5044 1004
rect 5164 996 5172 1004
rect 5676 996 5684 1004
rect 6188 996 6196 1004
rect 4620 976 4628 984
rect 4812 976 4820 984
rect 4908 976 4916 984
rect 5836 976 5844 984
rect 6252 980 6260 988
rect 172 956 180 964
rect 300 956 308 964
rect 428 956 436 964
rect 684 956 692 964
rect 716 956 724 964
rect 1292 956 1300 964
rect 1388 956 1396 964
rect 1484 956 1492 964
rect 1868 956 1876 964
rect 1996 956 2004 964
rect 2220 956 2228 964
rect 2284 956 2292 964
rect 3372 956 3380 964
rect 3692 956 3700 964
rect 4268 956 4276 964
rect 4428 956 4436 964
rect 4460 956 4468 964
rect 5100 956 5108 964
rect 5132 956 5140 964
rect 5228 956 5236 964
rect 5324 956 5332 964
rect 5420 956 5428 964
rect 5516 956 5524 964
rect 5612 956 5620 964
rect 5996 956 6004 964
rect 6252 956 6260 960
rect 6252 952 6260 956
rect 140 936 148 944
rect 812 936 820 944
rect 1036 936 1044 944
rect 684 916 692 924
rect 2444 936 2452 944
rect 2732 936 2740 944
rect 2764 936 2772 944
rect 2828 936 2836 944
rect 2988 936 2996 944
rect 3052 936 3060 944
rect 3084 936 3092 944
rect 1772 916 1780 924
rect 1804 916 1812 924
rect 2060 916 2068 924
rect 2620 916 2628 924
rect 2668 916 2676 924
rect 2796 916 2804 924
rect 3660 936 3668 944
rect 4012 936 4020 944
rect 4908 936 4916 944
rect 5004 936 5012 944
rect 5292 936 5300 944
rect 5484 940 5492 948
rect 5932 936 5940 944
rect 6124 936 6132 944
rect 652 896 660 904
rect 812 896 820 904
rect 908 896 916 904
rect 1548 896 1556 904
rect 1644 896 1652 904
rect 1868 896 1876 904
rect 2252 896 2260 904
rect 2316 896 2324 904
rect 2540 896 2548 904
rect 2572 896 2580 904
rect 2924 896 2932 904
rect 3212 896 3220 904
rect 3500 916 3508 924
rect 3532 916 3540 924
rect 3564 916 3572 924
rect 4140 916 4148 924
rect 4460 916 4468 924
rect 4620 916 4628 924
rect 3884 896 3892 904
rect 4108 896 4116 904
rect 4332 896 4340 904
rect 4588 896 4596 904
rect 4876 916 4884 924
rect 5084 916 5092 924
rect 5164 916 5172 924
rect 5484 912 5492 920
rect 4812 896 4820 904
rect 5004 896 5012 904
rect 5068 896 5076 904
rect 5228 896 5236 904
rect 5900 916 5908 924
rect 940 876 948 884
rect 1164 876 1172 884
rect 1260 876 1268 884
rect 1388 876 1396 884
rect 2860 876 2868 884
rect 3308 876 3316 884
rect 972 856 980 864
rect 1100 856 1108 864
rect 1196 856 1204 864
rect 2092 856 2100 864
rect 2252 856 2260 864
rect 2284 856 2292 864
rect 2444 856 2452 864
rect 2924 856 2932 864
rect 3532 856 3540 864
rect 3660 856 3668 864
rect 4300 876 4308 884
rect 4428 876 4436 884
rect 4556 876 4564 884
rect 4972 876 4980 884
rect 5100 876 5108 884
rect 5388 876 5396 884
rect 5932 896 5940 904
rect 6156 896 6164 904
rect 5900 876 5908 884
rect 4940 856 4948 864
rect 5356 856 5364 864
rect 5388 856 5396 864
rect 5676 856 5684 864
rect 5772 860 5780 868
rect 5996 856 6004 864
rect 6252 856 6260 864
rect 780 836 788 844
rect 1324 836 1332 844
rect 2348 836 2356 844
rect 2412 836 2420 844
rect 2636 836 2644 844
rect 3308 836 3316 844
rect 3340 836 3348 844
rect 3500 836 3508 844
rect 4108 836 4116 844
rect 5052 836 5060 844
rect 5772 832 5780 840
rect 5964 836 5972 844
rect 1068 816 1076 824
rect 2188 816 2196 824
rect 2348 816 2356 824
rect 1578 806 1585 814
rect 1585 806 1586 814
rect 1590 806 1595 814
rect 1595 806 1597 814
rect 1597 806 1598 814
rect 1602 806 1605 814
rect 1605 806 1607 814
rect 1607 806 1610 814
rect 1614 806 1615 814
rect 1615 806 1622 814
rect 1388 796 1396 804
rect 1420 796 1428 804
rect 460 776 468 784
rect 1068 776 1076 784
rect 1516 776 1524 784
rect 1676 796 1684 804
rect 1740 796 1748 804
rect 2060 796 2068 804
rect 2156 796 2164 804
rect 2300 796 2308 804
rect 2764 796 2772 804
rect 3052 796 3060 804
rect 4300 796 4308 804
rect 4332 816 4340 824
rect 4428 816 4436 824
rect 4588 816 4596 824
rect 5324 816 5332 824
rect 5420 816 5428 824
rect 4666 806 4673 814
rect 4673 806 4674 814
rect 4678 806 4683 814
rect 4683 806 4685 814
rect 4685 806 4686 814
rect 4690 806 4693 814
rect 4693 806 4695 814
rect 4695 806 4698 814
rect 4702 806 4703 814
rect 4703 806 4710 814
rect 4396 796 4404 804
rect 4748 796 4756 804
rect 4972 796 4980 804
rect 1900 776 1908 784
rect 2508 776 2516 784
rect 2988 776 2996 784
rect 4492 776 4500 784
rect 4940 776 4948 784
rect 5068 776 5076 784
rect 5260 776 5268 784
rect 1100 756 1108 764
rect 1452 756 1460 764
rect 1836 756 1844 764
rect 1868 756 1876 764
rect 2028 756 2036 764
rect 2124 756 2132 764
rect 1324 736 1332 744
rect 588 716 596 724
rect 812 716 820 724
rect 972 716 980 724
rect 940 696 948 704
rect 1964 736 1972 744
rect 2252 756 2260 764
rect 2284 756 2292 764
rect 2828 756 2836 764
rect 3340 756 3348 764
rect 5356 776 5364 784
rect 5932 776 5940 784
rect 5964 776 5972 784
rect 6060 776 6068 784
rect 6124 776 6132 784
rect 2188 736 2196 744
rect 2220 736 2228 744
rect 1868 716 1876 724
rect 2124 716 2132 724
rect 2156 716 2164 724
rect 2252 716 2260 724
rect 2316 736 2324 744
rect 3020 736 3028 744
rect 3308 736 3316 744
rect 3468 736 3476 744
rect 2572 716 2580 724
rect 2604 716 2612 724
rect 2636 716 2644 724
rect 2828 716 2836 724
rect 3276 716 3284 724
rect 5100 736 5108 744
rect 5484 736 5492 744
rect 6060 736 6068 744
rect 4332 716 4340 724
rect 4748 716 4756 724
rect 5004 716 5012 724
rect 5932 716 5940 724
rect 1132 700 1140 708
rect 1260 696 1268 704
rect 332 676 340 684
rect 908 676 916 684
rect 1004 676 1012 684
rect 1132 672 1140 680
rect 2444 696 2452 704
rect 2028 676 2036 684
rect 2188 676 2196 684
rect 2412 676 2420 684
rect 140 656 148 664
rect 1068 656 1076 664
rect 1260 656 1268 664
rect 1772 656 1780 664
rect 2060 656 2068 664
rect 556 636 564 644
rect 748 636 756 644
rect 1164 640 1172 648
rect 1740 636 1748 644
rect 2220 636 2228 644
rect 2668 676 2676 684
rect 2828 676 2836 684
rect 3436 696 3444 704
rect 3628 696 3636 704
rect 3980 696 3988 704
rect 4300 696 4308 704
rect 3308 676 3316 684
rect 4012 676 4020 684
rect 4588 676 4596 684
rect 4748 676 4756 684
rect 4812 676 4820 684
rect 5196 696 5204 704
rect 5260 696 5268 704
rect 5356 696 5364 704
rect 5484 696 5492 704
rect 5516 696 5524 704
rect 5308 676 5316 684
rect 5340 676 5348 684
rect 3084 656 3092 664
rect 3244 656 3252 664
rect 3756 656 3764 664
rect 2588 636 2596 644
rect 2956 636 2964 644
rect 3052 636 3060 644
rect 812 616 820 624
rect 940 616 948 624
rect 1132 616 1140 624
rect 1164 612 1172 620
rect 1836 616 1844 624
rect 1868 616 1876 624
rect 1996 616 2004 624
rect 2060 616 2068 624
rect 2124 616 2132 624
rect 2668 616 2676 624
rect 2700 616 2708 624
rect 2924 616 2932 624
rect 3244 616 3252 624
rect 3436 616 3444 624
rect 3114 606 3121 614
rect 3121 606 3122 614
rect 3126 606 3131 614
rect 3131 606 3133 614
rect 3133 606 3134 614
rect 3138 606 3141 614
rect 3141 606 3143 614
rect 3143 606 3146 614
rect 3150 606 3151 614
rect 3151 606 3158 614
rect 1452 596 1460 604
rect 364 556 372 564
rect 1516 576 1524 584
rect 1740 576 1748 584
rect 2252 596 2260 604
rect 2380 596 2388 604
rect 2412 596 2420 604
rect 2796 576 2804 584
rect 4332 616 4340 624
rect 4428 616 4436 624
rect 4460 616 4468 624
rect 5228 656 5236 664
rect 5292 656 5300 664
rect 5324 656 5332 664
rect 5996 676 6004 684
rect 6156 676 6164 684
rect 6252 696 6260 704
rect 6220 676 6228 684
rect 4780 636 4788 644
rect 4876 636 4884 644
rect 6252 636 6260 644
rect 4620 616 4628 624
rect 5004 616 5012 624
rect 5356 616 5364 624
rect 5388 616 5396 624
rect 5420 616 5428 624
rect 4972 596 4980 604
rect 5068 596 5076 604
rect 5228 596 5236 604
rect 5260 596 5268 604
rect 5516 596 5524 604
rect 3276 576 3284 584
rect 3628 576 3636 584
rect 3756 576 3764 584
rect 3788 576 3796 584
rect 3948 576 3956 584
rect 492 516 500 524
rect 684 516 692 524
rect 1100 536 1108 544
rect 1132 536 1140 544
rect 1324 536 1332 544
rect 1676 536 1684 544
rect 940 516 948 524
rect 1036 516 1044 524
rect 556 496 564 504
rect 1324 496 1332 504
rect 1484 496 1492 504
rect 1676 496 1684 504
rect 1804 516 1812 524
rect 2092 556 2100 564
rect 2764 556 2772 564
rect 3212 556 3220 564
rect 3244 556 3252 564
rect 3308 556 3316 564
rect 3660 556 3668 564
rect 3980 556 3988 564
rect 4108 556 4116 564
rect 4428 576 4436 584
rect 4460 576 4468 584
rect 4524 576 4532 584
rect 4812 576 4820 584
rect 4940 576 4948 584
rect 5164 576 5172 584
rect 6284 596 6292 604
rect 5996 576 6004 584
rect 4748 560 4756 568
rect 5100 556 5108 564
rect 5292 556 5300 564
rect 2028 536 2036 544
rect 1932 516 1940 524
rect 1964 516 1972 524
rect 2220 516 2228 524
rect 2412 516 2420 524
rect 2668 536 2676 544
rect 2956 536 2964 544
rect 3500 536 3508 544
rect 3532 536 3540 544
rect 3820 536 3828 544
rect 4012 536 4020 544
rect 4140 536 4148 544
rect 4204 536 4212 544
rect 4268 536 4276 544
rect 2732 516 2740 524
rect 4748 532 4756 540
rect 4812 536 4820 544
rect 5228 536 5236 544
rect 5260 536 5268 544
rect 5548 556 5556 564
rect 6252 556 6260 564
rect 5836 536 5844 544
rect 2860 516 2868 524
rect 2988 516 2996 524
rect 3340 516 3348 524
rect 3372 516 3380 524
rect 2156 496 2164 504
rect 2636 496 2644 504
rect 2764 496 2772 504
rect 2828 496 2836 504
rect 3020 496 3028 504
rect 3052 496 3060 504
rect 3500 496 3508 504
rect 3724 496 3732 504
rect 3788 516 3796 524
rect 3916 516 3924 524
rect 4300 516 4308 524
rect 4460 516 4468 524
rect 4492 516 4500 524
rect 4908 516 4916 524
rect 5004 516 5012 524
rect 5068 516 5076 524
rect 5132 516 5140 524
rect 5452 516 5460 524
rect 6092 516 6100 524
rect 12 476 20 484
rect 844 476 852 484
rect 1196 476 1204 484
rect 2540 476 2548 484
rect 2796 476 2804 484
rect 2892 476 2900 484
rect 3468 476 3476 484
rect 4236 496 4244 504
rect 4268 496 4276 504
rect 4556 496 4564 504
rect 4748 496 4756 504
rect 4876 496 4884 504
rect 5356 496 5364 504
rect 5868 496 5876 504
rect 4012 476 4020 484
rect 4428 476 4436 484
rect 5516 476 5524 484
rect 5612 476 5620 484
rect 2316 456 2324 464
rect 3276 456 3284 464
rect 4172 456 4180 464
rect 4972 456 4980 464
rect 5036 456 5044 464
rect 5324 456 5332 464
rect 5356 456 5364 464
rect 5420 456 5428 464
rect 5964 456 5972 464
rect 1932 436 1940 444
rect 2124 436 2132 444
rect 2476 436 2484 444
rect 3756 436 3764 444
rect 844 416 852 424
rect 1578 406 1585 414
rect 1585 406 1586 414
rect 1590 406 1595 414
rect 1595 406 1597 414
rect 1597 406 1598 414
rect 1602 406 1605 414
rect 1605 406 1607 414
rect 1607 406 1610 414
rect 1614 406 1615 414
rect 1615 406 1622 414
rect 588 396 596 404
rect 1324 396 1332 404
rect 1484 396 1492 404
rect 1772 396 1780 404
rect 1804 416 1812 424
rect 2156 416 2164 424
rect 2764 416 2772 424
rect 2924 416 2932 424
rect 3724 416 3732 424
rect 3852 436 3860 444
rect 3948 436 3956 444
rect 4364 436 4372 444
rect 4396 416 4404 424
rect 2412 396 2420 404
rect 2892 396 2900 404
rect 2956 396 2964 404
rect 2988 396 2996 404
rect 3020 396 3028 404
rect 3244 396 3252 404
rect 4012 396 4020 404
rect 4236 396 4244 404
rect 4492 396 4500 404
rect 4524 396 4532 404
rect 4556 396 4564 404
rect 4972 416 4980 424
rect 5356 416 5364 424
rect 5548 416 5556 424
rect 5772 416 5780 424
rect 4666 406 4673 414
rect 4673 406 4674 414
rect 4678 406 4683 414
rect 4683 406 4685 414
rect 4685 406 4686 414
rect 4690 406 4693 414
rect 4693 406 4695 414
rect 4695 406 4698 414
rect 4702 406 4703 414
rect 4703 406 4710 414
rect 4876 396 4884 404
rect 5036 396 5044 404
rect 5932 396 5940 404
rect 140 376 148 384
rect 1132 376 1140 384
rect 3596 376 3604 384
rect 3692 376 3700 384
rect 3724 376 3732 384
rect 1068 336 1076 344
rect 1932 356 1940 364
rect 1964 356 1972 364
rect 2412 356 2420 364
rect 2796 356 2804 364
rect 3756 356 3764 364
rect 3852 356 3860 364
rect 4044 356 4052 364
rect 4812 376 4820 384
rect 5228 376 5236 384
rect 5964 376 5972 384
rect 5772 356 5780 364
rect 5932 356 5940 364
rect 876 316 884 324
rect 1324 316 1332 324
rect 492 296 500 304
rect 1292 300 1300 308
rect 2508 336 2516 344
rect 2540 336 2548 344
rect 1900 296 1908 304
rect 1932 296 1940 304
rect 1996 296 2004 304
rect 2156 296 2164 304
rect 2636 316 2644 324
rect 2348 296 2356 304
rect 2412 296 2420 304
rect 2508 296 2516 304
rect 236 276 244 284
rect 716 276 724 284
rect 1260 276 1268 284
rect 1292 272 1300 280
rect 1356 276 1364 284
rect 1420 276 1428 284
rect 1484 276 1492 284
rect 1516 276 1524 284
rect 1708 276 1716 284
rect 1772 276 1780 284
rect 364 256 372 264
rect 1228 256 1236 264
rect 2604 276 2612 284
rect 2764 296 2772 304
rect 2828 336 2836 344
rect 2956 336 2964 344
rect 3212 336 3220 344
rect 3436 336 3444 344
rect 3564 336 3572 344
rect 3660 336 3668 344
rect 3692 336 3700 344
rect 4780 336 4788 344
rect 2860 316 2868 324
rect 3532 316 3540 324
rect 3628 316 3636 324
rect 3852 316 3860 324
rect 4236 316 4244 324
rect 4268 316 4276 324
rect 2924 296 2932 304
rect 2988 296 2996 304
rect 2652 276 2660 284
rect 2700 276 2708 284
rect 3324 276 3332 284
rect 3404 276 3412 284
rect 3436 276 3444 284
rect 3628 276 3636 284
rect 3724 296 3732 304
rect 3932 276 3940 284
rect 4108 276 4116 284
rect 4140 276 4148 284
rect 4204 296 4212 304
rect 4524 316 4532 324
rect 4556 316 4564 324
rect 4588 316 4596 324
rect 4620 316 4628 324
rect 4780 296 4788 304
rect 4396 276 4404 284
rect 4556 276 4564 284
rect 2988 256 2996 264
rect 3532 256 3540 264
rect 3660 256 3668 264
rect 3852 256 3860 264
rect 3884 256 3892 264
rect 4076 256 4084 264
rect 4588 256 4596 264
rect 5004 296 5012 304
rect 5100 296 5108 304
rect 5132 296 5140 304
rect 5356 316 5364 324
rect 5676 336 5684 344
rect 6156 356 6164 364
rect 6060 316 6068 324
rect 5164 276 5172 284
rect 5676 276 5684 284
rect 5772 276 5780 284
rect 5868 296 5876 304
rect 5964 296 5972 304
rect 4844 256 4852 264
rect 4940 256 4948 264
rect 5036 256 5044 264
rect 5420 256 5428 264
rect 5452 256 5460 264
rect 5932 256 5940 264
rect 972 236 980 244
rect 1324 236 1332 244
rect 1532 236 1540 244
rect 1964 236 1972 244
rect 2156 236 2164 244
rect 2828 236 2836 244
rect 2892 236 2900 244
rect 4236 236 4244 244
rect 876 216 884 224
rect 1676 216 1684 224
rect 1900 216 1908 224
rect 1356 196 1364 204
rect 1500 196 1508 204
rect 1740 196 1748 204
rect 1772 196 1780 204
rect 1820 196 1828 204
rect 2316 196 2324 204
rect 2380 216 2388 224
rect 2668 216 2676 224
rect 3052 216 3060 224
rect 3114 206 3121 214
rect 3121 206 3122 214
rect 3126 206 3131 214
rect 3131 206 3133 214
rect 3133 206 3134 214
rect 3138 206 3141 214
rect 3141 206 3143 214
rect 3143 206 3146 214
rect 3150 206 3151 214
rect 3151 206 3158 214
rect 2796 196 2804 204
rect 2908 196 2916 204
rect 3244 196 3252 204
rect 3564 216 3572 224
rect 3596 216 3604 224
rect 3724 216 3732 224
rect 4492 236 4500 244
rect 4812 236 4820 244
rect 3756 196 3764 204
rect 4524 196 4532 204
rect 332 176 340 184
rect 780 176 788 184
rect 1964 176 1972 184
rect 2028 176 2036 184
rect 844 156 852 164
rect 1068 156 1076 164
rect 1260 156 1268 164
rect 1356 156 1364 164
rect 2092 176 2100 184
rect 3276 176 3284 184
rect 2060 136 2068 144
rect 2156 136 2164 144
rect 2828 156 2836 164
rect 2956 156 2964 164
rect 3324 156 3332 164
rect 3500 156 3508 164
rect 3532 156 3540 164
rect 4108 176 4116 184
rect 4332 156 4340 164
rect 5036 176 5044 184
rect 5276 196 5284 204
rect 5420 196 5428 204
rect 6156 196 6164 204
rect 5356 176 5364 184
rect 5644 176 5652 184
rect 4460 156 4468 164
rect 4876 156 4884 164
rect 5004 156 5012 164
rect 5132 156 5140 164
rect 5196 156 5204 164
rect 5900 176 5908 184
rect 5932 176 5940 184
rect 5804 156 5812 164
rect 6252 156 6260 164
rect 2316 136 2324 144
rect 3692 136 3700 144
rect 3724 136 3732 144
rect 3820 136 3828 144
rect 4300 136 4308 144
rect 5036 136 5044 144
rect 5580 136 5588 144
rect 5996 136 6004 144
rect 6156 136 6164 144
rect 492 116 500 124
rect 812 116 820 124
rect 972 116 980 124
rect 1164 116 1172 124
rect 1260 116 1268 124
rect 1516 116 1524 124
rect 1900 116 1908 124
rect 1964 116 1972 124
rect 2140 116 2148 124
rect 2220 116 2228 124
rect 2540 116 2548 124
rect 940 96 948 104
rect 1292 96 1300 104
rect 2060 96 2068 104
rect 2668 116 2676 124
rect 2732 96 2740 104
rect 3020 116 3028 124
rect 3052 116 3060 124
rect 3212 96 3220 104
rect 3340 96 3348 104
rect 3532 116 3540 124
rect 3564 116 3572 124
rect 3756 116 3764 124
rect 4396 116 4404 124
rect 4812 116 4820 124
rect 5292 116 5300 124
rect 5324 116 5332 124
rect 5388 116 5396 124
rect 5708 116 5716 124
rect 5740 116 5748 124
rect 6092 116 6100 124
rect 6188 116 6196 124
rect 3884 96 3892 104
rect 3980 96 3988 104
rect 4076 96 4084 104
rect 4108 96 4116 104
rect 5068 96 5076 104
rect 5676 96 5684 104
rect 6028 96 6036 104
rect 2492 76 2500 84
rect 2556 76 2564 84
rect 1548 56 1556 64
rect 2796 76 2804 84
rect 2828 76 2836 84
rect 4044 76 4052 84
rect 4508 76 4516 84
rect 4956 76 4964 84
rect 5196 76 5204 84
rect 5420 76 5428 84
rect 5932 76 5940 84
rect 3084 56 3092 64
rect 236 36 244 44
rect 2604 36 2612 44
rect 2828 36 2836 44
rect 3436 56 3444 64
rect 3660 56 3668 64
rect 4364 56 4372 64
rect 4428 56 4436 64
rect 4556 56 4564 64
rect 5004 56 5012 64
rect 5036 56 5044 64
rect 5452 56 5460 64
rect 5740 56 5748 64
rect 4012 36 4020 44
rect 2124 16 2132 24
rect 2700 16 2708 24
rect 4188 36 4196 44
rect 5260 36 5268 44
rect 5292 36 5300 44
rect 4140 16 4148 24
rect 5356 16 5364 24
rect 5388 16 5396 24
rect 5484 16 5492 24
rect 5740 16 5748 24
rect 6124 16 6132 24
rect 1578 6 1585 14
rect 1585 6 1586 14
rect 1590 6 1595 14
rect 1595 6 1597 14
rect 1597 6 1598 14
rect 1602 6 1605 14
rect 1605 6 1607 14
rect 1607 6 1610 14
rect 1614 6 1615 14
rect 1615 6 1622 14
rect 4666 6 4673 14
rect 4673 6 4674 14
rect 4678 6 4683 14
rect 4683 6 4685 14
rect 4685 6 4686 14
rect 4690 6 4693 14
rect 4693 6 4695 14
rect 4695 6 4698 14
rect 4702 6 4703 14
rect 4703 6 4710 14
<< metal4 >>
rect 522 4604 534 4606
rect 522 4596 524 4604
rect 532 4596 534 4604
rect 202 4544 214 4546
rect 202 4536 204 4544
rect 212 4536 214 4544
rect 138 4124 150 4126
rect 138 4116 140 4124
rect 148 4116 150 4124
rect 138 3864 150 4116
rect 202 4124 214 4536
rect 458 4524 470 4526
rect 458 4516 460 4524
rect 468 4516 470 4524
rect 202 4116 204 4124
rect 212 4116 214 4124
rect 202 4104 214 4116
rect 202 4096 204 4104
rect 212 4096 214 4104
rect 202 3924 214 4096
rect 202 3916 204 3924
rect 212 3916 214 3924
rect 138 3856 140 3864
rect 148 3856 150 3864
rect 138 3854 150 3856
rect 170 3904 182 3906
rect 170 3896 172 3904
rect 180 3896 182 3904
rect 138 3744 150 3746
rect 138 3736 140 3744
rect 148 3736 150 3744
rect 138 3644 150 3736
rect 138 3636 140 3644
rect 148 3636 150 3644
rect 138 3634 150 3636
rect 138 3604 150 3606
rect 138 3596 140 3604
rect 148 3596 150 3604
rect 10 3244 22 3246
rect 10 3236 12 3244
rect 20 3236 22 3244
rect 10 2524 22 3236
rect 138 3204 150 3596
rect 138 3196 140 3204
rect 148 3196 150 3204
rect 138 3194 150 3196
rect 138 3164 150 3166
rect 138 3156 140 3164
rect 148 3156 150 3164
rect 10 2516 12 2524
rect 20 2516 22 2524
rect 10 2514 22 2516
rect 106 2584 118 2586
rect 106 2576 108 2584
rect 116 2576 118 2584
rect 74 2384 86 2386
rect 74 2376 76 2384
rect 84 2376 86 2384
rect 10 2304 22 2306
rect 10 2296 12 2304
rect 20 2296 22 2304
rect 10 1104 22 2296
rect 74 1764 86 2376
rect 106 1904 118 2576
rect 138 2544 150 3156
rect 170 2764 182 3896
rect 170 2756 172 2764
rect 180 2756 182 2764
rect 170 2754 182 2756
rect 202 3864 214 3916
rect 202 3856 204 3864
rect 212 3856 214 3864
rect 202 3744 214 3856
rect 202 3736 204 3744
rect 212 3736 214 3744
rect 202 3704 214 3736
rect 202 3696 204 3704
rect 212 3696 214 3704
rect 202 3524 214 3696
rect 234 4364 246 4366
rect 234 4356 236 4364
rect 244 4356 246 4364
rect 234 3884 246 4356
rect 362 4184 374 4186
rect 362 4176 364 4184
rect 372 4176 374 4184
rect 362 4164 374 4176
rect 362 4156 364 4164
rect 372 4156 374 4164
rect 330 4104 342 4106
rect 330 4096 332 4104
rect 340 4096 342 4104
rect 330 3924 342 4096
rect 330 3916 332 3924
rect 340 3916 342 3924
rect 330 3914 342 3916
rect 234 3876 236 3884
rect 244 3876 246 3884
rect 234 3704 246 3876
rect 234 3696 236 3704
rect 244 3696 246 3704
rect 234 3694 246 3696
rect 266 3804 278 3806
rect 266 3796 268 3804
rect 276 3796 278 3804
rect 202 3516 204 3524
rect 212 3516 214 3524
rect 202 3084 214 3516
rect 234 3624 246 3626
rect 234 3616 236 3624
rect 244 3616 246 3624
rect 234 3104 246 3616
rect 266 3544 278 3796
rect 266 3536 268 3544
rect 276 3536 278 3544
rect 266 3534 278 3536
rect 298 3764 310 3766
rect 298 3756 300 3764
rect 308 3756 310 3764
rect 266 3504 278 3506
rect 266 3496 268 3504
rect 276 3496 278 3504
rect 266 3224 278 3496
rect 266 3216 268 3224
rect 276 3216 278 3224
rect 266 3214 278 3216
rect 234 3096 236 3104
rect 244 3096 246 3104
rect 234 3094 246 3096
rect 202 3076 204 3084
rect 212 3076 214 3084
rect 202 2564 214 3076
rect 202 2556 204 2564
rect 212 2556 214 2564
rect 202 2554 214 2556
rect 234 2824 246 2826
rect 234 2816 236 2824
rect 244 2816 246 2824
rect 138 2536 140 2544
rect 148 2536 150 2544
rect 138 2534 150 2536
rect 106 1896 108 1904
rect 116 1896 118 1904
rect 106 1894 118 1896
rect 170 2124 182 2126
rect 170 2116 172 2124
rect 180 2116 182 2124
rect 170 1864 182 2116
rect 170 1856 172 1864
rect 180 1856 182 1864
rect 170 1854 182 1856
rect 74 1756 76 1764
rect 84 1756 86 1764
rect 74 1754 86 1756
rect 234 1504 246 2816
rect 298 2544 310 3756
rect 362 3724 374 4156
rect 458 4084 470 4516
rect 458 4076 460 4084
rect 468 4076 470 4084
rect 458 4074 470 4076
rect 522 3924 534 4596
rect 746 4584 758 4586
rect 746 4576 748 4584
rect 756 4576 758 4584
rect 714 4524 726 4526
rect 714 4516 716 4524
rect 724 4516 726 4524
rect 522 3916 524 3924
rect 532 3916 534 3924
rect 522 3914 534 3916
rect 682 4144 694 4146
rect 682 4136 684 4144
rect 692 4136 694 4144
rect 554 3904 566 3906
rect 554 3896 556 3904
rect 564 3896 566 3904
rect 522 3884 534 3886
rect 522 3876 524 3884
rect 532 3876 534 3884
rect 362 3716 364 3724
rect 372 3716 374 3724
rect 362 3714 374 3716
rect 394 3804 406 3806
rect 394 3796 396 3804
rect 404 3796 406 3804
rect 394 3744 406 3796
rect 394 3736 396 3744
rect 404 3736 406 3744
rect 394 3524 406 3736
rect 426 3804 486 3806
rect 426 3796 476 3804
rect 484 3796 486 3804
rect 426 3794 486 3796
rect 426 3664 438 3794
rect 426 3656 428 3664
rect 436 3656 438 3664
rect 426 3654 438 3656
rect 458 3744 470 3746
rect 458 3736 460 3744
rect 468 3736 470 3744
rect 458 3664 470 3736
rect 458 3656 460 3664
rect 468 3656 470 3664
rect 458 3654 470 3656
rect 394 3516 396 3524
rect 404 3516 406 3524
rect 394 3514 406 3516
rect 490 3404 502 3406
rect 490 3396 492 3404
rect 500 3396 502 3404
rect 426 3224 438 3226
rect 426 3216 428 3224
rect 436 3216 438 3224
rect 330 3104 342 3106
rect 330 3096 332 3104
rect 340 3096 342 3104
rect 330 2964 342 3096
rect 330 2956 332 2964
rect 340 2956 342 2964
rect 330 2954 342 2956
rect 394 2924 406 2926
rect 394 2916 396 2924
rect 404 2916 406 2924
rect 362 2744 374 2746
rect 362 2736 364 2744
rect 372 2736 374 2744
rect 362 2684 374 2736
rect 362 2676 364 2684
rect 372 2676 374 2684
rect 362 2674 374 2676
rect 298 2536 300 2544
rect 308 2536 310 2544
rect 298 2534 310 2536
rect 394 2224 406 2916
rect 426 2704 438 3216
rect 426 2696 428 2704
rect 436 2696 438 2704
rect 426 2694 438 2696
rect 458 3124 470 3126
rect 458 3116 460 3124
rect 468 3116 470 3124
rect 458 2884 470 3116
rect 490 3024 502 3396
rect 490 3016 492 3024
rect 500 3016 502 3024
rect 490 3014 502 3016
rect 522 3384 534 3876
rect 554 3704 566 3896
rect 554 3696 556 3704
rect 564 3696 566 3704
rect 554 3694 566 3696
rect 618 3724 630 3726
rect 618 3716 620 3724
rect 628 3716 630 3724
rect 522 3376 524 3384
rect 532 3376 534 3384
rect 458 2876 460 2884
rect 468 2876 470 2884
rect 458 2664 470 2876
rect 490 2924 502 2926
rect 490 2916 492 2924
rect 500 2916 502 2924
rect 490 2804 502 2916
rect 490 2796 492 2804
rect 500 2796 502 2804
rect 490 2794 502 2796
rect 458 2656 460 2664
rect 468 2656 470 2664
rect 458 2624 470 2656
rect 458 2616 460 2624
rect 468 2616 470 2624
rect 458 2614 470 2616
rect 490 2684 502 2686
rect 490 2676 492 2684
rect 500 2676 502 2684
rect 458 2564 470 2566
rect 458 2556 460 2564
rect 468 2556 470 2564
rect 458 2404 470 2556
rect 490 2484 502 2676
rect 490 2476 492 2484
rect 500 2476 502 2484
rect 490 2474 502 2476
rect 522 2684 534 3376
rect 522 2676 524 2684
rect 532 2676 534 2684
rect 522 2544 534 2676
rect 522 2536 524 2544
rect 532 2536 534 2544
rect 458 2396 460 2404
rect 468 2396 470 2404
rect 458 2394 470 2396
rect 426 2344 438 2346
rect 426 2336 428 2344
rect 436 2336 438 2344
rect 426 2264 438 2336
rect 522 2304 534 2536
rect 522 2296 524 2304
rect 532 2296 534 2304
rect 522 2294 534 2296
rect 554 3544 566 3546
rect 554 3536 556 3544
rect 564 3536 566 3544
rect 554 3284 566 3536
rect 554 3276 556 3284
rect 564 3276 566 3284
rect 554 3144 566 3276
rect 586 3524 598 3526
rect 586 3516 588 3524
rect 596 3516 598 3524
rect 586 3364 598 3516
rect 618 3484 630 3716
rect 618 3476 620 3484
rect 628 3476 630 3484
rect 618 3474 630 3476
rect 650 3524 662 3526
rect 650 3516 652 3524
rect 660 3516 662 3524
rect 586 3356 588 3364
rect 596 3356 598 3364
rect 586 3164 598 3356
rect 586 3156 588 3164
rect 596 3156 598 3164
rect 586 3154 598 3156
rect 618 3324 630 3326
rect 618 3316 620 3324
rect 628 3316 630 3324
rect 554 3136 556 3144
rect 564 3136 566 3144
rect 554 2744 566 3136
rect 586 3124 598 3126
rect 586 3116 588 3124
rect 596 3116 598 3124
rect 586 3084 598 3116
rect 586 3076 588 3084
rect 596 3076 598 3084
rect 586 3074 598 3076
rect 618 3104 630 3316
rect 618 3096 620 3104
rect 628 3096 630 3104
rect 554 2736 556 2744
rect 564 2736 566 2744
rect 554 2504 566 2736
rect 554 2496 556 2504
rect 564 2496 566 2504
rect 426 2256 428 2264
rect 436 2256 438 2264
rect 426 2254 438 2256
rect 394 2216 396 2224
rect 404 2216 406 2224
rect 394 2214 406 2216
rect 426 2204 438 2206
rect 426 2196 428 2204
rect 436 2196 438 2204
rect 394 2124 406 2126
rect 394 2116 396 2124
rect 404 2116 406 2124
rect 362 2104 374 2106
rect 362 2096 364 2104
rect 372 2096 374 2104
rect 362 1904 374 2096
rect 394 1964 406 2116
rect 394 1956 396 1964
rect 404 1956 406 1964
rect 394 1954 406 1956
rect 362 1896 364 1904
rect 372 1896 374 1904
rect 362 1894 374 1896
rect 426 1524 438 2196
rect 490 2184 502 2186
rect 490 2176 492 2184
rect 500 2176 502 2184
rect 490 2024 502 2176
rect 490 2016 492 2024
rect 500 2016 502 2024
rect 490 2014 502 2016
rect 554 2084 566 2496
rect 586 3004 598 3006
rect 586 2996 588 3004
rect 596 2996 598 3004
rect 586 2144 598 2996
rect 586 2136 588 2144
rect 596 2136 598 2144
rect 586 2134 598 2136
rect 618 2704 630 3096
rect 650 2824 662 3516
rect 682 2984 694 4136
rect 714 3464 726 4516
rect 714 3456 716 3464
rect 724 3456 726 3464
rect 714 3004 726 3456
rect 714 2996 716 3004
rect 724 2996 726 3004
rect 714 2994 726 2996
rect 682 2976 684 2984
rect 692 2976 694 2984
rect 682 2974 694 2976
rect 650 2816 652 2824
rect 660 2816 662 2824
rect 650 2814 662 2816
rect 618 2696 620 2704
rect 628 2696 630 2704
rect 618 2544 630 2696
rect 682 2724 710 2726
rect 682 2716 700 2724
rect 708 2716 710 2724
rect 682 2714 710 2716
rect 682 2686 694 2714
rect 650 2674 694 2686
rect 650 2664 662 2674
rect 650 2656 652 2664
rect 660 2656 662 2664
rect 650 2654 662 2656
rect 714 2664 726 2666
rect 714 2656 716 2664
rect 724 2656 726 2664
rect 682 2624 694 2626
rect 682 2616 684 2624
rect 692 2616 694 2624
rect 618 2536 620 2544
rect 628 2536 630 2544
rect 618 2124 630 2536
rect 650 2544 662 2546
rect 650 2536 652 2544
rect 660 2536 662 2544
rect 650 2204 662 2536
rect 682 2464 694 2616
rect 714 2604 726 2656
rect 714 2596 716 2604
rect 724 2596 726 2604
rect 714 2594 726 2596
rect 682 2456 684 2464
rect 692 2456 694 2464
rect 682 2454 694 2456
rect 714 2564 726 2566
rect 714 2556 716 2564
rect 724 2556 726 2564
rect 714 2464 726 2556
rect 746 2484 758 4576
rect 1130 4544 1142 4546
rect 1130 4536 1132 4544
rect 1140 4536 1142 4544
rect 1098 4524 1110 4526
rect 1098 4516 1100 4524
rect 1108 4516 1110 4524
rect 1002 4324 1014 4326
rect 1002 4316 1004 4324
rect 1012 4316 1014 4324
rect 810 4244 822 4246
rect 810 4236 812 4244
rect 820 4236 822 4244
rect 810 3824 822 4236
rect 874 4244 886 4246
rect 874 4236 876 4244
rect 884 4236 886 4244
rect 874 4164 886 4236
rect 874 4156 876 4164
rect 884 4156 886 4164
rect 874 4154 886 4156
rect 970 4184 982 4186
rect 970 4176 972 4184
rect 980 4176 982 4184
rect 970 3864 982 4176
rect 1002 4104 1014 4316
rect 1034 4264 1046 4266
rect 1034 4256 1036 4264
rect 1044 4256 1046 4264
rect 1034 4144 1046 4256
rect 1034 4136 1036 4144
rect 1044 4136 1046 4144
rect 1034 4134 1046 4136
rect 1002 4096 1004 4104
rect 1012 4096 1014 4104
rect 1002 4094 1014 4096
rect 970 3856 972 3864
rect 980 3856 982 3864
rect 970 3854 982 3856
rect 1066 3864 1078 3866
rect 1066 3856 1068 3864
rect 1076 3856 1078 3864
rect 810 3816 812 3824
rect 820 3816 822 3824
rect 810 3814 822 3816
rect 1002 3844 1014 3846
rect 1002 3836 1004 3844
rect 1012 3836 1014 3844
rect 938 3804 950 3806
rect 938 3796 940 3804
rect 948 3796 950 3804
rect 906 3764 918 3766
rect 906 3756 908 3764
rect 916 3756 918 3764
rect 810 3584 822 3586
rect 810 3576 812 3584
rect 820 3576 822 3584
rect 810 3264 822 3576
rect 842 3564 854 3566
rect 842 3556 844 3564
rect 852 3556 854 3564
rect 842 3364 854 3556
rect 906 3524 918 3756
rect 906 3516 908 3524
rect 916 3516 918 3524
rect 906 3514 918 3516
rect 938 3404 950 3796
rect 938 3396 940 3404
rect 948 3396 950 3404
rect 938 3394 950 3396
rect 970 3644 982 3646
rect 970 3636 972 3644
rect 980 3636 982 3644
rect 842 3356 844 3364
rect 852 3356 854 3364
rect 842 3354 854 3356
rect 874 3384 886 3386
rect 874 3376 876 3384
rect 884 3376 886 3384
rect 810 3256 812 3264
rect 820 3256 822 3264
rect 810 3254 822 3256
rect 842 3184 854 3186
rect 842 3176 844 3184
rect 852 3176 854 3184
rect 778 3064 790 3066
rect 778 3056 780 3064
rect 788 3056 790 3064
rect 778 2964 790 3056
rect 842 3024 854 3176
rect 874 3084 886 3376
rect 906 3344 918 3346
rect 906 3336 908 3344
rect 916 3336 918 3344
rect 906 3104 918 3336
rect 906 3096 908 3104
rect 916 3096 918 3104
rect 906 3094 918 3096
rect 938 3164 950 3166
rect 938 3156 940 3164
rect 948 3156 950 3164
rect 874 3076 876 3084
rect 884 3076 886 3084
rect 874 3074 886 3076
rect 842 3016 844 3024
rect 852 3016 854 3024
rect 842 3014 854 3016
rect 778 2956 780 2964
rect 788 2956 790 2964
rect 778 2954 790 2956
rect 874 2944 886 2946
rect 874 2936 876 2944
rect 884 2936 886 2944
rect 842 2824 854 2826
rect 842 2816 844 2824
rect 852 2816 854 2824
rect 842 2604 854 2816
rect 842 2596 844 2604
rect 852 2596 854 2604
rect 842 2594 854 2596
rect 746 2476 748 2484
rect 756 2476 758 2484
rect 746 2474 758 2476
rect 810 2524 822 2526
rect 810 2516 812 2524
rect 820 2516 822 2524
rect 714 2456 716 2464
rect 724 2456 726 2464
rect 714 2454 726 2456
rect 682 2424 694 2426
rect 682 2416 684 2424
rect 692 2416 694 2424
rect 682 2406 694 2416
rect 682 2394 790 2406
rect 778 2364 790 2394
rect 778 2356 780 2364
rect 788 2356 790 2364
rect 778 2354 790 2356
rect 650 2196 652 2204
rect 660 2196 662 2204
rect 650 2194 662 2196
rect 682 2344 694 2346
rect 682 2336 684 2344
rect 692 2336 694 2344
rect 618 2116 620 2124
rect 628 2116 630 2124
rect 554 2076 556 2084
rect 564 2076 566 2084
rect 490 1964 502 1966
rect 490 1956 492 1964
rect 500 1956 502 1964
rect 426 1516 428 1524
rect 436 1516 438 1524
rect 426 1514 438 1516
rect 458 1684 470 1686
rect 458 1676 460 1684
rect 468 1676 470 1684
rect 234 1496 236 1504
rect 244 1496 246 1504
rect 234 1494 246 1496
rect 362 1484 374 1486
rect 362 1476 364 1484
rect 372 1476 374 1484
rect 266 1344 278 1346
rect 266 1336 268 1344
rect 276 1336 278 1344
rect 170 1324 182 1326
rect 170 1316 172 1324
rect 180 1316 182 1324
rect 10 1096 12 1104
rect 20 1096 22 1104
rect 10 484 22 1096
rect 74 1184 86 1186
rect 74 1176 76 1184
rect 84 1176 86 1184
rect 74 1024 86 1176
rect 74 1016 76 1024
rect 84 1016 86 1024
rect 74 1014 86 1016
rect 170 1124 182 1316
rect 170 1116 172 1124
rect 180 1116 182 1124
rect 170 964 182 1116
rect 266 1104 278 1336
rect 266 1096 268 1104
rect 276 1096 278 1104
rect 266 984 278 1096
rect 266 976 268 984
rect 276 976 278 984
rect 266 974 278 976
rect 298 1344 310 1346
rect 298 1336 300 1344
rect 308 1336 310 1344
rect 298 1064 310 1336
rect 298 1056 300 1064
rect 308 1056 310 1064
rect 170 956 172 964
rect 180 956 182 964
rect 170 954 182 956
rect 298 964 310 1056
rect 298 956 300 964
rect 308 956 310 964
rect 298 954 310 956
rect 10 476 12 484
rect 20 476 22 484
rect 10 474 22 476
rect 138 944 150 946
rect 138 936 140 944
rect 148 936 150 944
rect 138 664 150 936
rect 138 656 140 664
rect 148 656 150 664
rect 138 384 150 656
rect 138 376 140 384
rect 148 376 150 384
rect 138 374 150 376
rect 330 684 342 686
rect 330 676 332 684
rect 340 676 342 684
rect 234 284 246 286
rect 234 276 236 284
rect 244 276 246 284
rect 234 44 246 276
rect 330 184 342 676
rect 362 564 374 1476
rect 426 1004 438 1006
rect 426 996 428 1004
rect 436 996 438 1004
rect 426 964 438 996
rect 426 956 428 964
rect 436 956 438 964
rect 426 954 438 956
rect 458 784 470 1676
rect 458 776 460 784
rect 468 776 470 784
rect 458 774 470 776
rect 490 1564 502 1956
rect 490 1556 492 1564
rect 500 1556 502 1564
rect 362 556 364 564
rect 372 556 374 564
rect 362 264 374 556
rect 362 256 364 264
rect 372 256 374 264
rect 362 254 374 256
rect 490 524 502 1556
rect 554 1944 566 2076
rect 554 1936 556 1944
rect 564 1936 566 1944
rect 522 1504 534 1506
rect 522 1496 524 1504
rect 532 1496 534 1504
rect 522 1084 534 1496
rect 554 1504 566 1936
rect 586 2084 598 2086
rect 586 2076 588 2084
rect 596 2076 598 2084
rect 586 1704 598 2076
rect 618 1924 630 2116
rect 650 2164 662 2166
rect 650 2156 652 2164
rect 660 2156 662 2164
rect 650 2124 662 2156
rect 650 2116 652 2124
rect 660 2116 662 2124
rect 650 2114 662 2116
rect 618 1916 620 1924
rect 628 1916 630 1924
rect 618 1914 630 1916
rect 650 1944 662 1946
rect 650 1936 652 1944
rect 660 1936 662 1944
rect 650 1886 662 1936
rect 618 1874 662 1886
rect 618 1724 630 1874
rect 618 1716 620 1724
rect 628 1716 630 1724
rect 618 1714 630 1716
rect 586 1696 588 1704
rect 596 1696 598 1704
rect 586 1694 598 1696
rect 554 1496 556 1504
rect 564 1496 566 1504
rect 554 1494 566 1496
rect 522 1076 524 1084
rect 532 1076 534 1084
rect 522 1074 534 1076
rect 650 1064 662 1066
rect 650 1056 652 1064
rect 660 1056 662 1064
rect 650 904 662 1056
rect 682 964 694 2336
rect 778 2324 790 2326
rect 778 2316 780 2324
rect 788 2316 790 2324
rect 778 2244 790 2316
rect 778 2236 780 2244
rect 788 2236 790 2244
rect 778 2234 790 2236
rect 746 2204 758 2206
rect 746 2196 748 2204
rect 756 2196 758 2204
rect 714 1504 726 1506
rect 714 1496 716 1504
rect 724 1496 726 1504
rect 714 1324 726 1496
rect 746 1424 758 2196
rect 810 1744 822 2516
rect 842 2384 854 2386
rect 842 2376 844 2384
rect 852 2376 854 2384
rect 842 2224 854 2376
rect 842 2216 844 2224
rect 852 2216 854 2224
rect 842 2214 854 2216
rect 810 1736 812 1744
rect 820 1736 822 1744
rect 810 1524 822 1736
rect 810 1516 812 1524
rect 820 1516 822 1524
rect 746 1416 748 1424
rect 756 1416 758 1424
rect 746 1414 758 1416
rect 778 1504 790 1506
rect 778 1496 780 1504
rect 788 1496 790 1504
rect 714 1316 716 1324
rect 724 1316 726 1324
rect 714 1314 726 1316
rect 746 1164 758 1166
rect 746 1156 748 1164
rect 756 1156 758 1164
rect 714 1144 726 1146
rect 714 1136 716 1144
rect 724 1136 726 1144
rect 714 1004 726 1136
rect 714 996 716 1004
rect 724 996 726 1004
rect 714 994 726 996
rect 682 956 684 964
rect 692 956 694 964
rect 682 954 694 956
rect 714 964 726 966
rect 714 956 716 964
rect 724 956 726 964
rect 650 896 652 904
rect 660 896 662 904
rect 650 894 662 896
rect 682 924 694 926
rect 682 916 684 924
rect 692 916 694 924
rect 586 724 598 726
rect 586 716 588 724
rect 596 716 598 724
rect 490 516 492 524
rect 500 516 502 524
rect 490 304 502 516
rect 554 644 566 646
rect 554 636 556 644
rect 564 636 566 644
rect 554 504 566 636
rect 554 496 556 504
rect 564 496 566 504
rect 554 494 566 496
rect 586 404 598 716
rect 682 524 694 916
rect 682 516 684 524
rect 692 516 694 524
rect 682 514 694 516
rect 586 396 588 404
rect 596 396 598 404
rect 586 394 598 396
rect 490 296 492 304
rect 500 296 502 304
rect 330 176 332 184
rect 340 176 342 184
rect 330 174 342 176
rect 490 124 502 296
rect 714 284 726 956
rect 746 644 758 1156
rect 778 1064 790 1496
rect 810 1464 822 1516
rect 810 1456 812 1464
rect 820 1456 822 1464
rect 810 1454 822 1456
rect 842 2164 854 2166
rect 842 2156 844 2164
rect 852 2156 854 2164
rect 842 1844 854 2156
rect 874 1864 886 2936
rect 906 2904 918 2906
rect 906 2896 908 2904
rect 916 2896 918 2904
rect 906 2804 918 2896
rect 906 2796 908 2804
rect 916 2796 918 2804
rect 906 2024 918 2796
rect 906 2016 908 2024
rect 916 2016 918 2024
rect 906 2014 918 2016
rect 938 2764 950 3156
rect 970 3104 982 3636
rect 1002 3344 1014 3836
rect 1002 3336 1004 3344
rect 1012 3336 1014 3344
rect 1002 3334 1014 3336
rect 1034 3664 1046 3666
rect 1034 3656 1036 3664
rect 1044 3656 1046 3664
rect 1034 3344 1046 3656
rect 1034 3336 1036 3344
rect 1044 3336 1046 3344
rect 970 3096 972 3104
rect 980 3096 982 3104
rect 970 3094 982 3096
rect 1002 3244 1014 3246
rect 1002 3236 1004 3244
rect 1012 3236 1014 3244
rect 938 2756 940 2764
rect 948 2756 950 2764
rect 938 2024 950 2756
rect 970 3064 982 3066
rect 970 3056 972 3064
rect 980 3056 982 3064
rect 970 2564 982 3056
rect 1002 2944 1014 3236
rect 1034 3184 1046 3336
rect 1066 3244 1078 3856
rect 1098 3404 1110 4516
rect 1130 3964 1142 4536
rect 1576 4414 1624 4640
rect 1706 4624 1718 4626
rect 1706 4616 1708 4624
rect 1716 4616 1718 4624
rect 1706 4484 1718 4616
rect 2410 4624 2422 4626
rect 2410 4616 2412 4624
rect 2420 4616 2422 4624
rect 2058 4604 2070 4606
rect 2058 4596 2060 4604
rect 2068 4596 2070 4604
rect 1706 4476 1708 4484
rect 1716 4476 1718 4484
rect 1706 4474 1718 4476
rect 1802 4544 1814 4546
rect 1802 4536 1804 4544
rect 1812 4536 1814 4544
rect 1576 4406 1578 4414
rect 1586 4406 1590 4414
rect 1598 4406 1602 4414
rect 1610 4406 1614 4414
rect 1622 4406 1624 4414
rect 1258 4384 1270 4386
rect 1258 4376 1260 4384
rect 1268 4376 1270 4384
rect 1226 4124 1238 4126
rect 1226 4116 1228 4124
rect 1236 4116 1238 4124
rect 1226 4064 1238 4116
rect 1258 4124 1270 4376
rect 1514 4364 1526 4366
rect 1514 4356 1516 4364
rect 1524 4356 1526 4364
rect 1418 4264 1430 4266
rect 1418 4256 1420 4264
rect 1428 4256 1430 4264
rect 1386 4224 1398 4226
rect 1386 4216 1388 4224
rect 1396 4216 1398 4224
rect 1386 4206 1398 4216
rect 1258 4116 1260 4124
rect 1268 4116 1270 4124
rect 1258 4114 1270 4116
rect 1322 4194 1398 4206
rect 1226 4056 1228 4064
rect 1236 4056 1238 4064
rect 1226 4054 1238 4056
rect 1322 4064 1334 4194
rect 1322 4056 1324 4064
rect 1332 4056 1334 4064
rect 1322 4054 1334 4056
rect 1354 4144 1366 4146
rect 1354 4136 1356 4144
rect 1364 4136 1366 4144
rect 1354 4064 1366 4136
rect 1418 4144 1430 4256
rect 1418 4136 1420 4144
rect 1428 4136 1430 4144
rect 1418 4134 1430 4136
rect 1354 4056 1356 4064
rect 1364 4056 1366 4064
rect 1354 4054 1366 4056
rect 1290 4044 1302 4046
rect 1290 4036 1292 4044
rect 1300 4036 1302 4044
rect 1226 4024 1238 4026
rect 1226 4016 1228 4024
rect 1236 4016 1238 4024
rect 1194 3984 1206 3986
rect 1194 3976 1196 3984
rect 1204 3976 1206 3984
rect 1130 3956 1132 3964
rect 1140 3956 1142 3964
rect 1130 3954 1142 3956
rect 1162 3964 1174 3966
rect 1162 3956 1164 3964
rect 1172 3956 1174 3964
rect 1130 3764 1142 3766
rect 1130 3756 1132 3764
rect 1140 3756 1142 3764
rect 1130 3704 1142 3756
rect 1130 3696 1132 3704
rect 1140 3696 1142 3704
rect 1130 3694 1142 3696
rect 1098 3396 1100 3404
rect 1108 3396 1110 3404
rect 1098 3394 1110 3396
rect 1130 3604 1142 3606
rect 1130 3596 1132 3604
rect 1140 3596 1142 3604
rect 1130 3384 1142 3596
rect 1162 3584 1174 3956
rect 1194 3864 1206 3976
rect 1194 3856 1196 3864
rect 1204 3856 1206 3864
rect 1194 3854 1206 3856
rect 1226 3844 1238 4016
rect 1226 3836 1228 3844
rect 1236 3836 1238 3844
rect 1226 3834 1238 3836
rect 1258 3924 1270 3926
rect 1258 3916 1260 3924
rect 1268 3916 1270 3924
rect 1258 3844 1270 3916
rect 1258 3836 1260 3844
rect 1268 3836 1270 3844
rect 1258 3834 1270 3836
rect 1162 3576 1164 3584
rect 1172 3576 1174 3584
rect 1162 3574 1174 3576
rect 1194 3764 1206 3766
rect 1194 3756 1196 3764
rect 1204 3756 1206 3764
rect 1194 3564 1206 3756
rect 1194 3556 1196 3564
rect 1204 3556 1206 3564
rect 1194 3554 1206 3556
rect 1258 3524 1270 3526
rect 1258 3516 1260 3524
rect 1268 3516 1270 3524
rect 1130 3376 1132 3384
rect 1140 3376 1142 3384
rect 1130 3374 1142 3376
rect 1162 3464 1174 3466
rect 1162 3456 1164 3464
rect 1172 3456 1174 3464
rect 1066 3236 1068 3244
rect 1076 3236 1078 3244
rect 1066 3234 1078 3236
rect 1162 3324 1174 3456
rect 1258 3424 1270 3516
rect 1258 3416 1260 3424
rect 1268 3416 1270 3424
rect 1258 3414 1270 3416
rect 1162 3316 1164 3324
rect 1172 3316 1174 3324
rect 1034 3176 1036 3184
rect 1044 3176 1046 3184
rect 1034 3174 1046 3176
rect 1066 3184 1078 3186
rect 1066 3176 1068 3184
rect 1076 3176 1078 3184
rect 1002 2936 1004 2944
rect 1012 2936 1014 2944
rect 1002 2934 1014 2936
rect 1034 3104 1046 3106
rect 1034 3096 1036 3104
rect 1044 3096 1046 3104
rect 1034 2924 1046 3096
rect 1066 2944 1078 3176
rect 1162 2964 1174 3316
rect 1194 3404 1206 3406
rect 1194 3396 1196 3404
rect 1204 3396 1206 3404
rect 1194 3224 1206 3396
rect 1194 3216 1196 3224
rect 1204 3216 1206 3224
rect 1194 3214 1206 3216
rect 1226 3384 1238 3386
rect 1226 3376 1228 3384
rect 1236 3376 1238 3384
rect 1226 3204 1238 3376
rect 1226 3196 1228 3204
rect 1236 3196 1238 3204
rect 1226 3194 1238 3196
rect 1258 3384 1270 3386
rect 1258 3376 1260 3384
rect 1268 3376 1270 3384
rect 1258 3204 1270 3376
rect 1258 3196 1260 3204
rect 1268 3196 1270 3204
rect 1258 3194 1270 3196
rect 1290 3184 1302 4036
rect 1514 4044 1526 4356
rect 1514 4036 1516 4044
rect 1524 4036 1526 4044
rect 1514 4034 1526 4036
rect 1482 4024 1494 4026
rect 1482 4016 1484 4024
rect 1492 4016 1494 4024
rect 1386 3984 1398 3986
rect 1386 3976 1388 3984
rect 1396 3976 1398 3984
rect 1386 3724 1398 3976
rect 1450 3984 1462 3986
rect 1450 3976 1452 3984
rect 1460 3976 1462 3984
rect 1450 3944 1462 3976
rect 1450 3936 1452 3944
rect 1460 3936 1462 3944
rect 1450 3934 1462 3936
rect 1482 3924 1494 4016
rect 1576 4014 1624 4406
rect 1770 4404 1782 4406
rect 1770 4396 1772 4404
rect 1780 4396 1782 4404
rect 1738 4344 1750 4346
rect 1738 4336 1740 4344
rect 1748 4336 1750 4344
rect 1706 4244 1718 4246
rect 1706 4236 1708 4244
rect 1716 4236 1718 4244
rect 1658 4164 1686 4166
rect 1658 4156 1660 4164
rect 1668 4156 1686 4164
rect 1658 4154 1686 4156
rect 1674 4104 1686 4154
rect 1674 4096 1676 4104
rect 1684 4096 1686 4104
rect 1674 4094 1686 4096
rect 1706 4044 1718 4236
rect 1706 4036 1708 4044
rect 1716 4036 1718 4044
rect 1706 4034 1718 4036
rect 1576 4006 1578 4014
rect 1586 4006 1590 4014
rect 1598 4006 1602 4014
rect 1610 4006 1614 4014
rect 1622 4006 1624 4014
rect 1482 3916 1484 3924
rect 1492 3916 1494 3924
rect 1482 3914 1494 3916
rect 1514 4004 1526 4006
rect 1514 3996 1516 4004
rect 1524 3996 1526 4004
rect 1514 3864 1526 3996
rect 1514 3856 1516 3864
rect 1524 3856 1526 3864
rect 1514 3854 1526 3856
rect 1546 3884 1558 3886
rect 1546 3876 1548 3884
rect 1556 3876 1558 3884
rect 1418 3804 1430 3806
rect 1418 3796 1420 3804
rect 1428 3796 1430 3804
rect 1418 3764 1430 3796
rect 1418 3756 1420 3764
rect 1428 3756 1430 3764
rect 1418 3754 1430 3756
rect 1386 3716 1388 3724
rect 1396 3716 1398 3724
rect 1386 3624 1398 3716
rect 1386 3616 1388 3624
rect 1396 3616 1398 3624
rect 1322 3524 1334 3526
rect 1322 3516 1324 3524
rect 1332 3516 1334 3524
rect 1322 3404 1334 3516
rect 1322 3396 1324 3404
rect 1332 3396 1334 3404
rect 1322 3394 1334 3396
rect 1354 3524 1366 3526
rect 1354 3516 1356 3524
rect 1364 3516 1366 3524
rect 1354 3484 1366 3516
rect 1386 3524 1398 3616
rect 1450 3724 1462 3726
rect 1450 3716 1452 3724
rect 1460 3716 1462 3724
rect 1386 3516 1388 3524
rect 1396 3516 1398 3524
rect 1386 3514 1398 3516
rect 1418 3524 1430 3526
rect 1418 3516 1420 3524
rect 1428 3516 1430 3524
rect 1354 3476 1356 3484
rect 1364 3476 1366 3484
rect 1290 3176 1292 3184
rect 1300 3176 1302 3184
rect 1210 3164 1238 3166
rect 1210 3156 1212 3164
rect 1220 3156 1238 3164
rect 1210 3154 1238 3156
rect 1226 3126 1238 3154
rect 1290 3144 1302 3176
rect 1322 3364 1334 3366
rect 1322 3356 1324 3364
rect 1332 3356 1334 3364
rect 1322 3164 1334 3356
rect 1322 3156 1324 3164
rect 1332 3156 1334 3164
rect 1322 3154 1334 3156
rect 1290 3136 1292 3144
rect 1300 3136 1302 3144
rect 1290 3134 1302 3136
rect 1194 3124 1206 3126
rect 1194 3116 1196 3124
rect 1204 3116 1206 3124
rect 1194 3084 1206 3116
rect 1226 3124 1254 3126
rect 1226 3116 1244 3124
rect 1252 3116 1254 3124
rect 1226 3114 1254 3116
rect 1194 3076 1196 3084
rect 1204 3076 1206 3084
rect 1194 3074 1206 3076
rect 1258 3104 1270 3106
rect 1258 3096 1260 3104
rect 1268 3096 1270 3104
rect 1162 2956 1164 2964
rect 1172 2956 1174 2964
rect 1162 2954 1174 2956
rect 1226 2984 1238 2986
rect 1226 2976 1228 2984
rect 1236 2976 1238 2984
rect 1066 2936 1068 2944
rect 1076 2936 1078 2944
rect 1066 2934 1078 2936
rect 1034 2916 1036 2924
rect 1044 2916 1046 2924
rect 1034 2914 1046 2916
rect 1130 2924 1142 2926
rect 1130 2916 1132 2924
rect 1140 2916 1142 2924
rect 1066 2884 1078 2886
rect 1066 2876 1068 2884
rect 1076 2876 1078 2884
rect 1002 2704 1014 2706
rect 1002 2696 1004 2704
rect 1012 2696 1014 2704
rect 1002 2604 1014 2696
rect 1002 2596 1004 2604
rect 1012 2596 1014 2604
rect 1002 2594 1014 2596
rect 1034 2684 1046 2686
rect 1034 2676 1036 2684
rect 1044 2676 1046 2684
rect 970 2556 972 2564
rect 980 2556 982 2564
rect 970 2284 982 2556
rect 970 2276 972 2284
rect 980 2276 982 2284
rect 970 2274 982 2276
rect 1002 2344 1014 2346
rect 1002 2336 1004 2344
rect 1012 2336 1014 2344
rect 1002 2164 1014 2336
rect 1002 2156 1004 2164
rect 1012 2156 1014 2164
rect 1002 2154 1014 2156
rect 938 2016 940 2024
rect 948 2016 950 2024
rect 874 1856 876 1864
rect 884 1856 886 1864
rect 874 1854 886 1856
rect 842 1836 844 1844
rect 852 1836 854 1844
rect 842 1424 854 1836
rect 906 1664 918 1666
rect 906 1656 908 1664
rect 916 1656 918 1664
rect 842 1416 844 1424
rect 852 1416 854 1424
rect 842 1414 854 1416
rect 874 1564 886 1566
rect 874 1556 876 1564
rect 884 1556 886 1564
rect 842 1384 854 1386
rect 842 1376 844 1384
rect 852 1376 854 1384
rect 810 1144 822 1146
rect 810 1136 812 1144
rect 820 1136 822 1144
rect 810 1086 822 1136
rect 842 1144 854 1376
rect 874 1344 886 1556
rect 906 1404 918 1656
rect 938 1544 950 2016
rect 1034 2144 1046 2676
rect 1066 2684 1078 2876
rect 1066 2676 1068 2684
rect 1076 2676 1078 2684
rect 1066 2674 1078 2676
rect 1098 2724 1110 2726
rect 1098 2716 1100 2724
rect 1108 2716 1110 2724
rect 1066 2624 1078 2626
rect 1066 2616 1068 2624
rect 1076 2616 1078 2624
rect 1066 2204 1078 2616
rect 1098 2504 1110 2716
rect 1098 2496 1100 2504
rect 1108 2496 1110 2504
rect 1098 2494 1110 2496
rect 1066 2196 1068 2204
rect 1076 2196 1078 2204
rect 1066 2194 1078 2196
rect 1034 2136 1036 2144
rect 1044 2136 1046 2144
rect 1034 1984 1046 2136
rect 1066 2084 1078 2086
rect 1066 2076 1068 2084
rect 1076 2076 1078 2084
rect 1066 2024 1078 2076
rect 1066 2016 1068 2024
rect 1076 2016 1078 2024
rect 1066 2014 1078 2016
rect 1098 2084 1110 2086
rect 1098 2076 1100 2084
rect 1108 2076 1110 2084
rect 1034 1976 1036 1984
rect 1044 1976 1046 1984
rect 1034 1974 1046 1976
rect 1066 1824 1078 1826
rect 1066 1816 1068 1824
rect 1076 1816 1078 1824
rect 1034 1704 1046 1706
rect 1034 1696 1036 1704
rect 1044 1696 1046 1704
rect 1002 1644 1014 1646
rect 1002 1636 1004 1644
rect 1012 1636 1014 1644
rect 938 1536 940 1544
rect 948 1536 950 1544
rect 938 1534 950 1536
rect 970 1604 982 1606
rect 970 1596 972 1604
rect 980 1596 982 1604
rect 906 1396 908 1404
rect 916 1396 918 1404
rect 906 1394 918 1396
rect 874 1336 876 1344
rect 884 1336 886 1344
rect 874 1334 886 1336
rect 938 1364 950 1366
rect 938 1356 940 1364
rect 948 1356 950 1364
rect 938 1184 950 1356
rect 970 1204 982 1596
rect 1002 1584 1014 1636
rect 1002 1576 1004 1584
rect 1012 1576 1014 1584
rect 1002 1574 1014 1576
rect 1002 1464 1014 1466
rect 1002 1456 1004 1464
rect 1012 1456 1014 1464
rect 1002 1424 1014 1456
rect 1002 1416 1004 1424
rect 1012 1416 1014 1424
rect 1002 1414 1014 1416
rect 970 1196 972 1204
rect 980 1196 982 1204
rect 970 1194 982 1196
rect 1002 1304 1014 1306
rect 1002 1296 1004 1304
rect 1012 1296 1014 1304
rect 1002 1204 1014 1296
rect 1034 1264 1046 1696
rect 1066 1704 1078 1816
rect 1098 1764 1110 2076
rect 1130 2004 1142 2916
rect 1162 2904 1174 2906
rect 1162 2896 1164 2904
rect 1172 2896 1174 2904
rect 1162 2724 1174 2896
rect 1226 2844 1238 2976
rect 1258 2924 1270 3096
rect 1322 3064 1334 3066
rect 1322 3056 1324 3064
rect 1332 3056 1334 3064
rect 1322 2944 1334 3056
rect 1354 3044 1366 3476
rect 1418 3384 1430 3516
rect 1418 3376 1420 3384
rect 1428 3376 1430 3384
rect 1418 3374 1430 3376
rect 1386 3304 1398 3306
rect 1386 3296 1388 3304
rect 1396 3296 1398 3304
rect 1386 3084 1398 3296
rect 1418 3204 1430 3206
rect 1418 3196 1420 3204
rect 1428 3196 1430 3204
rect 1418 3124 1430 3196
rect 1418 3116 1420 3124
rect 1428 3116 1430 3124
rect 1418 3114 1430 3116
rect 1386 3076 1388 3084
rect 1396 3076 1398 3084
rect 1386 3074 1398 3076
rect 1354 3036 1356 3044
rect 1364 3036 1366 3044
rect 1354 3034 1366 3036
rect 1450 3004 1462 3716
rect 1546 3724 1558 3876
rect 1546 3716 1548 3724
rect 1556 3716 1558 3724
rect 1546 3714 1558 3716
rect 1482 3704 1494 3706
rect 1482 3696 1484 3704
rect 1492 3696 1494 3704
rect 1482 3544 1494 3696
rect 1576 3614 1624 4006
rect 1706 3804 1718 3806
rect 1706 3796 1708 3804
rect 1716 3796 1718 3804
rect 1674 3704 1686 3706
rect 1674 3696 1676 3704
rect 1684 3696 1686 3704
rect 1674 3624 1686 3696
rect 1674 3616 1676 3624
rect 1684 3616 1686 3624
rect 1674 3614 1686 3616
rect 1576 3606 1578 3614
rect 1586 3606 1590 3614
rect 1598 3606 1602 3614
rect 1610 3606 1614 3614
rect 1622 3606 1624 3614
rect 1482 3536 1484 3544
rect 1492 3536 1494 3544
rect 1482 3484 1494 3536
rect 1546 3544 1558 3546
rect 1546 3536 1548 3544
rect 1556 3536 1558 3544
rect 1482 3476 1484 3484
rect 1492 3476 1494 3484
rect 1482 3474 1494 3476
rect 1514 3504 1526 3506
rect 1514 3496 1516 3504
rect 1524 3496 1526 3504
rect 1514 3324 1526 3496
rect 1514 3316 1516 3324
rect 1524 3316 1526 3324
rect 1514 3314 1526 3316
rect 1546 3284 1558 3536
rect 1546 3276 1548 3284
rect 1556 3276 1558 3284
rect 1546 3274 1558 3276
rect 1514 3224 1526 3226
rect 1514 3216 1516 3224
rect 1524 3216 1526 3224
rect 1450 2996 1452 3004
rect 1460 2996 1462 3004
rect 1322 2936 1324 2944
rect 1332 2936 1334 2944
rect 1322 2934 1334 2936
rect 1418 2984 1430 2986
rect 1418 2976 1420 2984
rect 1428 2976 1430 2984
rect 1418 2944 1430 2976
rect 1450 2984 1462 2996
rect 1450 2976 1452 2984
rect 1460 2976 1462 2984
rect 1450 2974 1462 2976
rect 1482 3104 1494 3106
rect 1482 3096 1484 3104
rect 1492 3096 1494 3104
rect 1418 2936 1420 2944
rect 1428 2936 1430 2944
rect 1418 2934 1430 2936
rect 1258 2916 1260 2924
rect 1268 2916 1270 2924
rect 1258 2914 1270 2916
rect 1482 2904 1494 3096
rect 1514 3004 1526 3216
rect 1576 3214 1624 3606
rect 1706 3564 1718 3796
rect 1738 3804 1750 4336
rect 1738 3796 1740 3804
rect 1748 3796 1750 3804
rect 1738 3794 1750 3796
rect 1770 4304 1782 4396
rect 1770 4296 1772 4304
rect 1780 4296 1782 4304
rect 1770 3788 1782 4296
rect 1802 4064 1814 4536
rect 1898 4504 1910 4506
rect 1898 4496 1900 4504
rect 1908 4496 1910 4504
rect 1802 4056 1804 4064
rect 1812 4056 1814 4064
rect 1802 4054 1814 4056
rect 1834 4084 1846 4086
rect 1834 4076 1836 4084
rect 1844 4076 1846 4084
rect 1834 4046 1846 4076
rect 1818 4044 1846 4046
rect 1818 4036 1820 4044
rect 1828 4036 1846 4044
rect 1818 4034 1846 4036
rect 1866 4084 1878 4086
rect 1866 4076 1868 4084
rect 1876 4076 1878 4084
rect 1866 3984 1878 4076
rect 1866 3976 1868 3984
rect 1876 3976 1878 3984
rect 1866 3974 1878 3976
rect 1866 3924 1878 3926
rect 1866 3916 1868 3924
rect 1876 3916 1878 3924
rect 1802 3884 1814 3886
rect 1802 3876 1804 3884
rect 1812 3876 1814 3884
rect 1802 3844 1814 3876
rect 1802 3836 1804 3844
rect 1812 3836 1814 3844
rect 1802 3834 1814 3836
rect 1834 3884 1846 3886
rect 1834 3876 1836 3884
rect 1844 3876 1846 3884
rect 1770 3780 1772 3788
rect 1780 3780 1782 3788
rect 1770 3774 1782 3780
rect 1770 3760 1782 3766
rect 1770 3752 1772 3760
rect 1780 3752 1782 3760
rect 1706 3556 1708 3564
rect 1716 3556 1718 3564
rect 1706 3554 1718 3556
rect 1738 3704 1750 3706
rect 1738 3696 1740 3704
rect 1748 3696 1750 3704
rect 1706 3484 1718 3486
rect 1706 3476 1708 3484
rect 1716 3476 1718 3484
rect 1576 3206 1578 3214
rect 1586 3206 1590 3214
rect 1598 3206 1602 3214
rect 1610 3206 1614 3214
rect 1622 3206 1624 3214
rect 1530 3084 1558 3086
rect 1530 3076 1532 3084
rect 1540 3076 1558 3084
rect 1530 3074 1558 3076
rect 1514 2996 1516 3004
rect 1524 2996 1526 3004
rect 1514 2994 1526 2996
rect 1482 2896 1484 2904
rect 1492 2896 1494 2904
rect 1482 2894 1494 2896
rect 1546 2904 1558 3074
rect 1546 2896 1548 2904
rect 1556 2896 1558 2904
rect 1546 2894 1558 2896
rect 1226 2836 1228 2844
rect 1236 2836 1238 2844
rect 1226 2834 1238 2836
rect 1290 2844 1302 2846
rect 1290 2836 1292 2844
rect 1300 2836 1302 2844
rect 1258 2824 1270 2826
rect 1258 2816 1260 2824
rect 1268 2816 1270 2824
rect 1226 2804 1238 2806
rect 1226 2796 1228 2804
rect 1236 2796 1238 2804
rect 1162 2716 1164 2724
rect 1172 2716 1174 2724
rect 1162 2714 1174 2716
rect 1194 2784 1206 2786
rect 1194 2776 1196 2784
rect 1204 2776 1206 2784
rect 1162 2684 1174 2686
rect 1162 2676 1164 2684
rect 1172 2676 1174 2684
rect 1162 2644 1174 2676
rect 1194 2664 1206 2776
rect 1226 2764 1238 2796
rect 1258 2784 1270 2816
rect 1258 2776 1260 2784
rect 1268 2776 1270 2784
rect 1258 2774 1270 2776
rect 1226 2756 1228 2764
rect 1236 2756 1238 2764
rect 1226 2754 1238 2756
rect 1194 2656 1196 2664
rect 1204 2656 1206 2664
rect 1194 2654 1206 2656
rect 1258 2744 1270 2746
rect 1258 2736 1260 2744
rect 1268 2736 1270 2744
rect 1258 2684 1270 2736
rect 1258 2676 1260 2684
rect 1268 2676 1270 2684
rect 1162 2636 1164 2644
rect 1172 2636 1174 2644
rect 1162 2624 1174 2636
rect 1162 2616 1164 2624
rect 1172 2616 1174 2624
rect 1162 2614 1174 2616
rect 1194 2524 1206 2526
rect 1194 2516 1196 2524
rect 1204 2516 1206 2524
rect 1130 1996 1132 2004
rect 1140 1996 1142 2004
rect 1130 1994 1142 1996
rect 1162 2484 1174 2486
rect 1162 2476 1164 2484
rect 1172 2476 1174 2484
rect 1098 1756 1100 1764
rect 1108 1756 1110 1764
rect 1098 1754 1110 1756
rect 1130 1884 1142 1886
rect 1130 1876 1132 1884
rect 1140 1876 1142 1884
rect 1066 1696 1068 1704
rect 1076 1696 1078 1704
rect 1066 1694 1078 1696
rect 1130 1664 1142 1876
rect 1162 1824 1174 2476
rect 1194 2124 1206 2516
rect 1194 2116 1196 2124
rect 1204 2116 1206 2124
rect 1194 2114 1206 2116
rect 1258 2144 1270 2676
rect 1290 2544 1302 2836
rect 1576 2814 1624 3206
rect 1674 3324 1686 3326
rect 1674 3316 1676 3324
rect 1684 3316 1686 3324
rect 1642 3144 1654 3146
rect 1642 3136 1644 3144
rect 1652 3136 1654 3144
rect 1642 3004 1654 3136
rect 1674 3124 1686 3316
rect 1706 3324 1718 3476
rect 1706 3316 1708 3324
rect 1716 3316 1718 3324
rect 1706 3314 1718 3316
rect 1674 3116 1676 3124
rect 1684 3116 1686 3124
rect 1674 3114 1686 3116
rect 1706 3264 1718 3266
rect 1706 3256 1708 3264
rect 1716 3256 1718 3264
rect 1706 3064 1718 3256
rect 1738 3264 1750 3696
rect 1770 3484 1782 3752
rect 1802 3724 1814 3726
rect 1802 3716 1804 3724
rect 1812 3716 1814 3724
rect 1802 3504 1814 3716
rect 1834 3644 1846 3876
rect 1834 3636 1836 3644
rect 1844 3636 1846 3644
rect 1834 3634 1846 3636
rect 1802 3496 1804 3504
rect 1812 3496 1814 3504
rect 1802 3494 1814 3496
rect 1834 3604 1846 3606
rect 1834 3596 1836 3604
rect 1844 3596 1846 3604
rect 1770 3476 1772 3484
rect 1780 3476 1782 3484
rect 1770 3474 1782 3476
rect 1834 3404 1846 3596
rect 1866 3604 1878 3916
rect 1898 3764 1910 4496
rect 1930 4484 1942 4486
rect 1930 4476 1932 4484
rect 1940 4476 1942 4484
rect 1930 4384 1942 4476
rect 1930 4376 1932 4384
rect 1940 4376 1942 4384
rect 1930 4374 1942 4376
rect 1962 4314 2038 4326
rect 1962 4284 1974 4314
rect 1962 4276 1964 4284
rect 1972 4276 1974 4284
rect 1962 4274 1974 4276
rect 1994 4284 2006 4286
rect 1994 4276 1996 4284
rect 2004 4276 2006 4284
rect 1962 4104 1974 4106
rect 1962 4096 1964 4104
rect 1972 4096 1974 4104
rect 1898 3756 1900 3764
rect 1908 3756 1910 3764
rect 1898 3754 1910 3756
rect 1930 4064 1942 4066
rect 1930 4056 1932 4064
rect 1940 4056 1942 4064
rect 1866 3596 1868 3604
rect 1876 3596 1878 3604
rect 1866 3594 1878 3596
rect 1898 3564 1910 3566
rect 1898 3556 1900 3564
rect 1908 3556 1910 3564
rect 1834 3396 1836 3404
rect 1844 3396 1846 3404
rect 1834 3394 1846 3396
rect 1866 3484 1878 3486
rect 1866 3476 1868 3484
rect 1876 3476 1878 3484
rect 1802 3324 1814 3326
rect 1802 3316 1804 3324
rect 1812 3316 1814 3324
rect 1738 3256 1740 3264
rect 1748 3256 1750 3264
rect 1738 3254 1750 3256
rect 1770 3264 1782 3266
rect 1770 3256 1772 3264
rect 1780 3256 1782 3264
rect 1770 3224 1782 3256
rect 1770 3216 1772 3224
rect 1780 3216 1782 3224
rect 1770 3214 1782 3216
rect 1770 3104 1782 3106
rect 1770 3096 1772 3104
rect 1780 3096 1782 3104
rect 1706 3056 1708 3064
rect 1716 3056 1718 3064
rect 1706 3054 1718 3056
rect 1738 3084 1750 3086
rect 1738 3076 1740 3084
rect 1748 3076 1750 3084
rect 1642 2996 1644 3004
rect 1652 2996 1654 3004
rect 1642 2994 1654 2996
rect 1674 3024 1686 3026
rect 1674 3016 1676 3024
rect 1684 3016 1686 3024
rect 1576 2806 1578 2814
rect 1586 2806 1590 2814
rect 1598 2806 1602 2814
rect 1610 2806 1614 2814
rect 1622 2806 1624 2814
rect 1290 2536 1292 2544
rect 1300 2536 1302 2544
rect 1290 2534 1302 2536
rect 1354 2804 1366 2806
rect 1354 2796 1356 2804
rect 1364 2796 1366 2804
rect 1354 2524 1366 2796
rect 1482 2804 1494 2806
rect 1482 2796 1484 2804
rect 1492 2796 1494 2804
rect 1450 2764 1462 2766
rect 1450 2756 1452 2764
rect 1460 2756 1462 2764
rect 1354 2516 1356 2524
rect 1364 2516 1366 2524
rect 1354 2514 1366 2516
rect 1386 2724 1398 2726
rect 1386 2716 1388 2724
rect 1396 2716 1398 2724
rect 1322 2504 1334 2506
rect 1322 2496 1324 2504
rect 1332 2496 1334 2504
rect 1258 2136 1260 2144
rect 1268 2136 1270 2144
rect 1226 2104 1238 2106
rect 1226 2096 1228 2104
rect 1236 2096 1238 2104
rect 1162 1816 1164 1824
rect 1172 1816 1174 1824
rect 1162 1814 1174 1816
rect 1194 2004 1206 2006
rect 1194 1996 1196 2004
rect 1204 1996 1206 2004
rect 1194 1704 1206 1996
rect 1226 1864 1238 2096
rect 1226 1856 1228 1864
rect 1236 1856 1238 1864
rect 1226 1854 1238 1856
rect 1194 1696 1196 1704
rect 1204 1696 1206 1704
rect 1194 1694 1206 1696
rect 1130 1656 1132 1664
rect 1140 1656 1142 1664
rect 1130 1654 1142 1656
rect 1258 1664 1270 2136
rect 1290 2344 1302 2346
rect 1290 2336 1292 2344
rect 1300 2336 1302 2344
rect 1290 1924 1302 2336
rect 1322 2064 1334 2496
rect 1386 2344 1398 2716
rect 1418 2664 1430 2666
rect 1418 2656 1420 2664
rect 1428 2656 1430 2664
rect 1418 2444 1430 2656
rect 1418 2436 1420 2444
rect 1428 2436 1430 2444
rect 1418 2434 1430 2436
rect 1450 2444 1462 2756
rect 1482 2644 1494 2796
rect 1482 2636 1484 2644
rect 1492 2636 1494 2644
rect 1482 2634 1494 2636
rect 1514 2784 1526 2786
rect 1514 2776 1516 2784
rect 1524 2776 1526 2784
rect 1514 2606 1526 2776
rect 1482 2594 1526 2606
rect 1482 2584 1494 2594
rect 1482 2576 1484 2584
rect 1492 2576 1494 2584
rect 1482 2574 1494 2576
rect 1514 2584 1526 2586
rect 1514 2576 1516 2584
rect 1524 2576 1526 2584
rect 1514 2566 1526 2576
rect 1514 2564 1558 2566
rect 1514 2556 1548 2564
rect 1556 2556 1558 2564
rect 1514 2554 1558 2556
rect 1450 2436 1452 2444
rect 1460 2436 1462 2444
rect 1450 2434 1462 2436
rect 1514 2484 1526 2486
rect 1514 2476 1516 2484
rect 1524 2476 1526 2484
rect 1514 2364 1526 2476
rect 1514 2356 1516 2364
rect 1524 2356 1526 2364
rect 1514 2354 1526 2356
rect 1576 2414 1624 2806
rect 1674 2704 1686 3016
rect 1738 2924 1750 3076
rect 1738 2916 1740 2924
rect 1748 2916 1750 2924
rect 1738 2914 1750 2916
rect 1738 2864 1750 2866
rect 1738 2856 1740 2864
rect 1748 2856 1750 2864
rect 1674 2696 1676 2704
rect 1684 2696 1686 2704
rect 1674 2694 1686 2696
rect 1706 2764 1718 2766
rect 1706 2756 1708 2764
rect 1716 2756 1718 2764
rect 1576 2406 1578 2414
rect 1586 2406 1590 2414
rect 1598 2406 1602 2414
rect 1610 2406 1614 2414
rect 1622 2406 1624 2414
rect 1386 2336 1388 2344
rect 1396 2336 1398 2344
rect 1386 2334 1398 2336
rect 1450 2344 1462 2346
rect 1450 2336 1452 2344
rect 1460 2336 1462 2344
rect 1354 2284 1366 2286
rect 1354 2276 1356 2284
rect 1364 2276 1366 2284
rect 1354 2166 1366 2276
rect 1418 2184 1430 2186
rect 1418 2176 1420 2184
rect 1428 2176 1430 2184
rect 1354 2154 1398 2166
rect 1386 2144 1398 2154
rect 1386 2136 1388 2144
rect 1396 2136 1398 2144
rect 1386 2134 1398 2136
rect 1322 2056 1324 2064
rect 1332 2056 1334 2064
rect 1322 2054 1334 2056
rect 1386 2084 1398 2086
rect 1386 2076 1388 2084
rect 1396 2076 1398 2084
rect 1386 2024 1398 2076
rect 1386 2016 1388 2024
rect 1396 2016 1398 2024
rect 1354 2004 1366 2006
rect 1354 1996 1356 2004
rect 1364 1996 1366 2004
rect 1290 1916 1292 1924
rect 1300 1916 1302 1924
rect 1290 1914 1302 1916
rect 1322 1924 1334 1926
rect 1322 1916 1324 1924
rect 1332 1916 1334 1924
rect 1290 1884 1302 1886
rect 1290 1876 1292 1884
rect 1300 1876 1302 1884
rect 1290 1824 1302 1876
rect 1290 1816 1292 1824
rect 1300 1816 1302 1824
rect 1290 1814 1302 1816
rect 1322 1824 1334 1916
rect 1322 1816 1324 1824
rect 1332 1816 1334 1824
rect 1322 1814 1334 1816
rect 1354 1824 1366 1996
rect 1354 1816 1356 1824
rect 1364 1816 1366 1824
rect 1354 1814 1366 1816
rect 1386 1964 1398 2016
rect 1418 2006 1430 2176
rect 1402 2004 1430 2006
rect 1402 1996 1404 2004
rect 1412 1996 1430 2004
rect 1402 1994 1430 1996
rect 1386 1956 1388 1964
rect 1396 1956 1398 1964
rect 1386 1824 1398 1956
rect 1418 1964 1430 1966
rect 1418 1956 1420 1964
rect 1428 1956 1430 1964
rect 1418 1844 1430 1956
rect 1418 1836 1420 1844
rect 1428 1836 1430 1844
rect 1418 1834 1430 1836
rect 1386 1816 1388 1824
rect 1396 1816 1398 1824
rect 1386 1814 1398 1816
rect 1258 1656 1260 1664
rect 1268 1656 1270 1664
rect 1258 1654 1270 1656
rect 1322 1724 1334 1726
rect 1322 1716 1324 1724
rect 1332 1716 1334 1724
rect 1066 1644 1078 1646
rect 1066 1636 1068 1644
rect 1076 1636 1078 1644
rect 1066 1304 1078 1636
rect 1098 1624 1110 1626
rect 1098 1616 1100 1624
rect 1108 1616 1110 1624
rect 1098 1544 1110 1616
rect 1098 1536 1100 1544
rect 1108 1536 1110 1544
rect 1098 1534 1110 1536
rect 1258 1624 1270 1626
rect 1258 1616 1260 1624
rect 1268 1616 1270 1624
rect 1130 1524 1142 1526
rect 1130 1516 1132 1524
rect 1140 1516 1142 1524
rect 1066 1296 1068 1304
rect 1076 1296 1078 1304
rect 1066 1294 1078 1296
rect 1098 1404 1110 1406
rect 1098 1396 1100 1404
rect 1108 1396 1110 1404
rect 1034 1256 1036 1264
rect 1044 1256 1046 1264
rect 1034 1254 1046 1256
rect 1002 1196 1004 1204
rect 1012 1196 1014 1204
rect 1002 1194 1014 1196
rect 938 1176 940 1184
rect 948 1176 950 1184
rect 938 1174 950 1176
rect 1066 1184 1078 1186
rect 1066 1176 1068 1184
rect 1076 1176 1078 1184
rect 842 1136 844 1144
rect 852 1136 854 1144
rect 842 1134 854 1136
rect 874 1154 982 1166
rect 874 1086 886 1154
rect 938 1124 950 1126
rect 938 1116 940 1124
rect 948 1116 950 1124
rect 810 1074 886 1086
rect 906 1104 918 1106
rect 906 1096 908 1104
rect 916 1096 918 1104
rect 778 1056 780 1064
rect 788 1056 790 1064
rect 778 1054 790 1056
rect 810 1034 886 1046
rect 810 1004 822 1034
rect 810 996 812 1004
rect 820 996 822 1004
rect 810 994 822 996
rect 842 1004 854 1006
rect 842 996 844 1004
rect 852 996 854 1004
rect 810 944 822 946
rect 810 936 812 944
rect 820 936 822 944
rect 810 904 822 936
rect 810 896 812 904
rect 820 896 822 904
rect 746 636 748 644
rect 756 636 758 644
rect 746 634 758 636
rect 778 844 790 846
rect 778 836 780 844
rect 788 836 790 844
rect 714 276 716 284
rect 724 276 726 284
rect 714 274 726 276
rect 778 184 790 836
rect 810 724 822 896
rect 810 716 812 724
rect 820 716 822 724
rect 810 714 822 716
rect 778 176 780 184
rect 788 176 790 184
rect 778 174 790 176
rect 810 624 822 626
rect 810 616 812 624
rect 820 616 822 624
rect 490 116 492 124
rect 500 116 502 124
rect 490 114 502 116
rect 810 124 822 616
rect 842 484 854 996
rect 874 1004 886 1034
rect 874 996 876 1004
rect 884 996 886 1004
rect 874 994 886 996
rect 906 904 918 1096
rect 906 896 908 904
rect 916 896 918 904
rect 906 684 918 896
rect 938 884 950 1116
rect 970 1124 982 1154
rect 970 1116 972 1124
rect 980 1116 982 1124
rect 970 1114 982 1116
rect 986 1004 1014 1006
rect 986 996 988 1004
rect 996 996 1014 1004
rect 986 994 1014 996
rect 938 876 940 884
rect 948 876 950 884
rect 938 874 950 876
rect 970 864 982 866
rect 970 856 972 864
rect 980 856 982 864
rect 970 724 982 856
rect 970 716 972 724
rect 980 716 982 724
rect 970 714 982 716
rect 906 676 908 684
rect 916 676 918 684
rect 906 674 918 676
rect 938 704 950 706
rect 938 696 940 704
rect 948 696 950 704
rect 938 624 950 696
rect 1002 684 1014 994
rect 1066 1004 1078 1176
rect 1098 1126 1110 1396
rect 1130 1184 1142 1516
rect 1226 1524 1238 1526
rect 1226 1516 1228 1524
rect 1236 1516 1238 1524
rect 1194 1464 1206 1466
rect 1194 1456 1196 1464
rect 1204 1456 1206 1464
rect 1162 1424 1174 1426
rect 1162 1416 1164 1424
rect 1172 1416 1174 1424
rect 1162 1324 1174 1416
rect 1162 1316 1164 1324
rect 1172 1316 1174 1324
rect 1162 1314 1174 1316
rect 1130 1176 1132 1184
rect 1140 1176 1142 1184
rect 1130 1174 1142 1176
rect 1162 1284 1174 1286
rect 1162 1276 1164 1284
rect 1172 1276 1174 1284
rect 1162 1184 1174 1276
rect 1162 1176 1164 1184
rect 1172 1176 1174 1184
rect 1162 1174 1174 1176
rect 1098 1114 1142 1126
rect 1066 996 1068 1004
rect 1076 996 1078 1004
rect 1002 676 1004 684
rect 1012 676 1014 684
rect 1002 674 1014 676
rect 1034 944 1046 946
rect 1034 936 1036 944
rect 1044 936 1046 944
rect 938 616 940 624
rect 948 616 950 624
rect 938 614 950 616
rect 842 476 844 484
rect 852 476 854 484
rect 842 474 854 476
rect 938 524 950 526
rect 938 516 940 524
rect 948 516 950 524
rect 842 424 854 426
rect 842 416 844 424
rect 852 416 854 424
rect 842 164 854 416
rect 874 324 886 326
rect 874 316 876 324
rect 884 316 886 324
rect 874 224 886 316
rect 874 216 876 224
rect 884 216 886 224
rect 874 214 886 216
rect 842 156 844 164
rect 852 156 854 164
rect 842 154 854 156
rect 810 116 812 124
rect 820 116 822 124
rect 810 114 822 116
rect 938 104 950 516
rect 1034 524 1046 936
rect 1066 824 1078 996
rect 1098 1084 1110 1086
rect 1098 1076 1100 1084
rect 1108 1076 1110 1084
rect 1098 864 1110 1076
rect 1130 984 1142 1114
rect 1130 976 1132 984
rect 1140 976 1142 984
rect 1130 974 1142 976
rect 1162 1004 1174 1006
rect 1162 996 1164 1004
rect 1172 996 1174 1004
rect 1162 926 1174 996
rect 1194 1004 1206 1456
rect 1226 1444 1238 1516
rect 1258 1484 1270 1616
rect 1258 1476 1260 1484
rect 1268 1476 1270 1484
rect 1258 1474 1270 1476
rect 1290 1524 1302 1526
rect 1290 1516 1292 1524
rect 1300 1516 1302 1524
rect 1226 1436 1228 1444
rect 1236 1436 1238 1444
rect 1226 1434 1238 1436
rect 1258 1444 1270 1446
rect 1258 1436 1260 1444
rect 1268 1436 1270 1444
rect 1194 996 1196 1004
rect 1204 996 1206 1004
rect 1194 994 1206 996
rect 1226 1384 1238 1386
rect 1226 1376 1228 1384
rect 1236 1376 1238 1384
rect 1098 856 1100 864
rect 1108 856 1110 864
rect 1098 854 1110 856
rect 1130 914 1174 926
rect 1066 816 1068 824
rect 1076 816 1078 824
rect 1066 814 1078 816
rect 1066 784 1078 786
rect 1066 776 1068 784
rect 1076 776 1078 784
rect 1066 664 1078 776
rect 1066 656 1068 664
rect 1076 656 1078 664
rect 1066 654 1078 656
rect 1098 764 1110 766
rect 1098 756 1100 764
rect 1108 756 1110 764
rect 1098 544 1110 756
rect 1130 708 1142 914
rect 1130 700 1132 708
rect 1140 700 1142 708
rect 1130 694 1142 700
rect 1162 884 1174 886
rect 1162 876 1164 884
rect 1172 876 1174 884
rect 1130 680 1142 686
rect 1130 672 1132 680
rect 1140 672 1142 680
rect 1130 624 1142 672
rect 1162 648 1174 876
rect 1162 640 1164 648
rect 1172 640 1174 648
rect 1162 634 1174 640
rect 1194 864 1206 866
rect 1194 856 1196 864
rect 1204 856 1206 864
rect 1130 616 1132 624
rect 1140 616 1142 624
rect 1130 614 1142 616
rect 1162 620 1174 626
rect 1162 612 1164 620
rect 1172 612 1174 620
rect 1098 536 1100 544
rect 1108 536 1110 544
rect 1098 534 1110 536
rect 1130 544 1142 546
rect 1130 536 1132 544
rect 1140 536 1142 544
rect 1034 516 1036 524
rect 1044 516 1046 524
rect 1034 514 1046 516
rect 1130 384 1142 536
rect 1130 376 1132 384
rect 1140 376 1142 384
rect 1130 374 1142 376
rect 1066 344 1078 346
rect 1066 336 1068 344
rect 1076 336 1078 344
rect 970 244 982 246
rect 970 236 972 244
rect 980 236 982 244
rect 970 124 982 236
rect 1066 164 1078 336
rect 1066 156 1068 164
rect 1076 156 1078 164
rect 1066 154 1078 156
rect 970 116 972 124
rect 980 116 982 124
rect 970 114 982 116
rect 1162 124 1174 612
rect 1194 484 1206 856
rect 1194 476 1196 484
rect 1204 476 1206 484
rect 1194 474 1206 476
rect 1226 264 1238 1376
rect 1258 1284 1270 1436
rect 1290 1324 1302 1516
rect 1290 1316 1292 1324
rect 1300 1316 1302 1324
rect 1290 1314 1302 1316
rect 1258 1276 1260 1284
rect 1268 1276 1270 1284
rect 1258 1274 1270 1276
rect 1290 1204 1302 1206
rect 1290 1196 1292 1204
rect 1300 1196 1302 1204
rect 1258 1104 1270 1106
rect 1258 1096 1260 1104
rect 1268 1096 1270 1104
rect 1258 884 1270 1096
rect 1290 964 1302 1196
rect 1290 956 1292 964
rect 1300 956 1302 964
rect 1290 954 1302 956
rect 1258 876 1260 884
rect 1268 876 1270 884
rect 1258 874 1270 876
rect 1322 844 1334 1716
rect 1418 1724 1430 1726
rect 1418 1716 1420 1724
rect 1428 1716 1430 1724
rect 1386 1664 1398 1666
rect 1386 1656 1388 1664
rect 1396 1656 1398 1664
rect 1354 1624 1366 1626
rect 1354 1616 1356 1624
rect 1364 1616 1366 1624
rect 1354 1584 1366 1616
rect 1354 1576 1356 1584
rect 1364 1576 1366 1584
rect 1354 1574 1366 1576
rect 1354 1424 1366 1426
rect 1354 1416 1356 1424
rect 1364 1416 1366 1424
rect 1354 1364 1366 1416
rect 1354 1356 1356 1364
rect 1364 1356 1366 1364
rect 1354 1354 1366 1356
rect 1386 1364 1398 1656
rect 1418 1464 1430 1716
rect 1450 1504 1462 2336
rect 1576 2014 1624 2406
rect 1674 2484 1686 2486
rect 1674 2476 1676 2484
rect 1684 2476 1686 2484
rect 1642 2364 1654 2366
rect 1642 2356 1644 2364
rect 1652 2356 1654 2364
rect 1642 2324 1654 2356
rect 1642 2316 1644 2324
rect 1652 2316 1654 2324
rect 1642 2314 1654 2316
rect 1642 2144 1654 2146
rect 1642 2136 1644 2144
rect 1652 2136 1654 2144
rect 1642 2064 1654 2136
rect 1674 2144 1686 2476
rect 1706 2484 1718 2756
rect 1738 2744 1750 2856
rect 1770 2844 1782 3096
rect 1802 3084 1814 3316
rect 1834 3324 1846 3326
rect 1834 3316 1836 3324
rect 1844 3316 1846 3324
rect 1834 3104 1846 3316
rect 1834 3096 1836 3104
rect 1844 3096 1846 3104
rect 1834 3094 1846 3096
rect 1802 3076 1804 3084
rect 1812 3076 1814 3084
rect 1802 3074 1814 3076
rect 1834 3064 1846 3066
rect 1834 3056 1836 3064
rect 1844 3056 1846 3064
rect 1834 2966 1846 3056
rect 1866 3004 1878 3476
rect 1898 3364 1910 3556
rect 1898 3356 1900 3364
rect 1908 3356 1910 3364
rect 1898 3354 1910 3356
rect 1930 3304 1942 4056
rect 1962 3544 1974 4096
rect 1994 4064 2006 4276
rect 2026 4284 2038 4314
rect 2026 4276 2028 4284
rect 2036 4276 2038 4284
rect 2026 4274 2038 4276
rect 1994 4056 1996 4064
rect 2004 4056 2006 4064
rect 1994 4054 2006 4056
rect 2026 4184 2038 4186
rect 2026 4176 2028 4184
rect 2036 4176 2038 4184
rect 2026 4024 2038 4176
rect 2058 4124 2070 4596
rect 2122 4604 2134 4606
rect 2122 4596 2124 4604
rect 2132 4596 2134 4604
rect 2058 4116 2060 4124
rect 2068 4116 2070 4124
rect 2058 4114 2070 4116
rect 2090 4224 2102 4226
rect 2090 4216 2092 4224
rect 2100 4216 2102 4224
rect 2026 4016 2028 4024
rect 2036 4016 2038 4024
rect 2026 4014 2038 4016
rect 2058 3984 2070 3986
rect 2058 3976 2060 3984
rect 2068 3976 2070 3984
rect 2026 3944 2038 3946
rect 2026 3936 2028 3944
rect 2036 3936 2038 3944
rect 1962 3536 1964 3544
rect 1972 3536 1974 3544
rect 1962 3534 1974 3536
rect 1994 3924 2006 3926
rect 1994 3916 1996 3924
rect 2004 3916 2006 3924
rect 1994 3544 2006 3916
rect 2026 3624 2038 3936
rect 2058 3904 2070 3976
rect 2058 3896 2060 3904
rect 2068 3896 2070 3904
rect 2058 3894 2070 3896
rect 2026 3616 2028 3624
rect 2036 3616 2038 3624
rect 2026 3614 2038 3616
rect 2058 3844 2070 3846
rect 2058 3836 2060 3844
rect 2068 3836 2070 3844
rect 1994 3536 1996 3544
rect 2004 3536 2006 3544
rect 1994 3534 2006 3536
rect 2026 3564 2038 3566
rect 2026 3556 2028 3564
rect 2036 3556 2038 3564
rect 1962 3464 1974 3466
rect 1962 3456 1964 3464
rect 1972 3456 1974 3464
rect 1962 3404 1974 3456
rect 1962 3396 1964 3404
rect 1972 3396 1974 3404
rect 1962 3394 1974 3396
rect 1994 3364 2006 3366
rect 1994 3356 1996 3364
rect 2004 3356 2006 3364
rect 1930 3296 1932 3304
rect 1940 3296 1942 3304
rect 1930 3294 1942 3296
rect 1962 3304 1974 3306
rect 1962 3296 1964 3304
rect 1972 3296 1974 3304
rect 1898 3244 1910 3246
rect 1898 3236 1900 3244
rect 1908 3236 1910 3244
rect 1898 3064 1910 3236
rect 1898 3056 1900 3064
rect 1908 3056 1910 3064
rect 1898 3054 1910 3056
rect 1866 2996 1868 3004
rect 1876 2996 1878 3004
rect 1866 2994 1878 2996
rect 1898 3024 1910 3026
rect 1898 3016 1900 3024
rect 1908 3016 1910 3024
rect 1802 2964 1814 2966
rect 1802 2956 1804 2964
rect 1812 2956 1814 2964
rect 1802 2864 1814 2956
rect 1834 2954 1878 2966
rect 1802 2856 1804 2864
rect 1812 2856 1814 2864
rect 1802 2854 1814 2856
rect 1834 2904 1846 2906
rect 1834 2896 1836 2904
rect 1844 2896 1846 2904
rect 1770 2836 1772 2844
rect 1780 2836 1782 2844
rect 1770 2834 1782 2836
rect 1738 2736 1740 2744
rect 1748 2736 1750 2744
rect 1738 2734 1750 2736
rect 1770 2784 1782 2786
rect 1770 2776 1772 2784
rect 1780 2776 1782 2784
rect 1770 2686 1782 2776
rect 1834 2704 1846 2896
rect 1866 2884 1878 2954
rect 1866 2876 1868 2884
rect 1876 2876 1878 2884
rect 1866 2874 1878 2876
rect 1834 2696 1836 2704
rect 1844 2696 1846 2704
rect 1834 2694 1846 2696
rect 1866 2844 1878 2846
rect 1866 2836 1868 2844
rect 1876 2836 1878 2844
rect 1754 2684 1782 2686
rect 1754 2676 1756 2684
rect 1764 2676 1782 2684
rect 1754 2674 1782 2676
rect 1866 2664 1878 2836
rect 1866 2656 1868 2664
rect 1876 2656 1878 2664
rect 1866 2654 1878 2656
rect 1706 2476 1708 2484
rect 1716 2476 1718 2484
rect 1706 2474 1718 2476
rect 1770 2644 1782 2646
rect 1770 2636 1772 2644
rect 1780 2636 1782 2644
rect 1738 2284 1750 2286
rect 1738 2276 1740 2284
rect 1748 2276 1750 2284
rect 1738 2184 1750 2276
rect 1738 2176 1740 2184
rect 1748 2176 1750 2184
rect 1674 2136 1676 2144
rect 1684 2136 1686 2144
rect 1674 2134 1686 2136
rect 1706 2164 1718 2166
rect 1706 2156 1708 2164
rect 1716 2156 1718 2164
rect 1706 2124 1718 2156
rect 1706 2116 1708 2124
rect 1716 2116 1718 2124
rect 1706 2114 1718 2116
rect 1738 2124 1750 2176
rect 1770 2164 1782 2636
rect 1834 2644 1846 2646
rect 1834 2636 1836 2644
rect 1844 2636 1846 2644
rect 1834 2404 1846 2636
rect 1834 2396 1836 2404
rect 1844 2396 1846 2404
rect 1834 2394 1846 2396
rect 1866 2624 1878 2626
rect 1866 2616 1868 2624
rect 1876 2616 1878 2624
rect 1866 2244 1878 2616
rect 1898 2446 1910 3016
rect 1930 3024 1942 3026
rect 1930 3016 1932 3024
rect 1940 3016 1942 3024
rect 1930 2544 1942 3016
rect 1962 2824 1974 3296
rect 1994 3064 2006 3356
rect 2026 3264 2038 3556
rect 2058 3304 2070 3836
rect 2090 3704 2102 4216
rect 2090 3696 2092 3704
rect 2100 3696 2102 3704
rect 2090 3694 2102 3696
rect 2058 3296 2060 3304
rect 2068 3296 2070 3304
rect 2058 3294 2070 3296
rect 2090 3444 2102 3446
rect 2090 3436 2092 3444
rect 2100 3436 2102 3444
rect 2090 3404 2102 3436
rect 2090 3396 2092 3404
rect 2100 3396 2102 3404
rect 2026 3256 2028 3264
rect 2036 3256 2038 3264
rect 2026 3254 2038 3256
rect 2090 3244 2102 3396
rect 2122 3324 2134 4596
rect 2314 4544 2326 4546
rect 2314 4536 2316 4544
rect 2324 4536 2326 4544
rect 2314 4364 2326 4536
rect 2314 4356 2316 4364
rect 2324 4356 2326 4364
rect 2314 4354 2326 4356
rect 2378 4444 2390 4446
rect 2378 4436 2380 4444
rect 2388 4436 2390 4444
rect 2186 4284 2342 4286
rect 2186 4276 2188 4284
rect 2196 4276 2332 4284
rect 2340 4276 2342 4284
rect 2186 4274 2342 4276
rect 2346 4184 2358 4186
rect 2346 4176 2348 4184
rect 2356 4176 2358 4184
rect 2186 4104 2198 4106
rect 2186 4096 2188 4104
rect 2196 4096 2198 4104
rect 2122 3316 2124 3324
rect 2132 3316 2134 3324
rect 2122 3314 2134 3316
rect 2154 4024 2166 4026
rect 2154 4016 2156 4024
rect 2164 4016 2166 4024
rect 2154 3924 2166 4016
rect 2154 3916 2156 3924
rect 2164 3916 2166 3924
rect 2154 3264 2166 3916
rect 2154 3256 2156 3264
rect 2164 3256 2166 3264
rect 2154 3254 2166 3256
rect 2186 3704 2198 4096
rect 2314 4044 2326 4046
rect 2314 4036 2316 4044
rect 2324 4036 2326 4044
rect 2314 3904 2326 4036
rect 2314 3896 2316 3904
rect 2324 3896 2326 3904
rect 2314 3894 2326 3896
rect 2186 3696 2188 3704
rect 2196 3696 2198 3704
rect 2186 3504 2198 3696
rect 2218 3804 2230 3806
rect 2218 3796 2220 3804
rect 2228 3796 2230 3804
rect 2218 3584 2230 3796
rect 2314 3724 2326 3726
rect 2314 3716 2316 3724
rect 2324 3716 2326 3724
rect 2282 3704 2294 3706
rect 2282 3696 2284 3704
rect 2292 3696 2294 3704
rect 2218 3576 2220 3584
rect 2228 3576 2230 3584
rect 2218 3574 2230 3576
rect 2250 3684 2262 3686
rect 2250 3676 2252 3684
rect 2260 3676 2262 3684
rect 2186 3496 2188 3504
rect 2196 3496 2198 3504
rect 2090 3236 2092 3244
rect 2100 3236 2102 3244
rect 2090 3234 2102 3236
rect 2122 3244 2134 3246
rect 2122 3236 2124 3244
rect 2132 3236 2134 3244
rect 2090 3184 2102 3186
rect 2090 3176 2092 3184
rect 2100 3176 2102 3184
rect 2058 3144 2070 3146
rect 2058 3136 2060 3144
rect 2068 3136 2070 3144
rect 1994 3056 1996 3064
rect 2004 3056 2006 3064
rect 1994 3054 2006 3056
rect 2026 3064 2038 3066
rect 2026 3056 2028 3064
rect 2036 3056 2038 3064
rect 1962 2816 1964 2824
rect 1972 2816 1974 2824
rect 1962 2744 1974 2816
rect 1994 2964 2006 2966
rect 1994 2956 1996 2964
rect 2004 2956 2006 2964
rect 1994 2804 2006 2956
rect 1994 2796 1996 2804
rect 2004 2796 2006 2804
rect 1994 2794 2006 2796
rect 1962 2736 1964 2744
rect 1972 2736 1974 2744
rect 1962 2734 1974 2736
rect 1994 2744 2006 2746
rect 1994 2736 1996 2744
rect 2004 2736 2006 2744
rect 1994 2704 2006 2736
rect 1994 2696 1996 2704
rect 2004 2696 2006 2704
rect 1994 2694 2006 2696
rect 1930 2536 1932 2544
rect 1940 2536 1942 2544
rect 1930 2534 1942 2536
rect 1962 2644 1974 2646
rect 1962 2636 1964 2644
rect 1972 2636 1974 2644
rect 1898 2434 1942 2446
rect 1866 2236 1868 2244
rect 1876 2236 1878 2244
rect 1770 2156 1772 2164
rect 1780 2156 1782 2164
rect 1770 2154 1782 2156
rect 1802 2224 1814 2226
rect 1802 2216 1804 2224
rect 1812 2216 1814 2224
rect 1738 2116 1740 2124
rect 1748 2116 1750 2124
rect 1738 2114 1750 2116
rect 1802 2124 1814 2216
rect 1866 2204 1878 2236
rect 1866 2196 1868 2204
rect 1876 2196 1878 2204
rect 1866 2194 1878 2196
rect 1802 2116 1804 2124
rect 1812 2116 1814 2124
rect 1802 2114 1814 2116
rect 1834 2184 1846 2186
rect 1834 2176 1836 2184
rect 1844 2176 1846 2184
rect 1802 2084 1814 2086
rect 1802 2076 1804 2084
rect 1812 2076 1814 2084
rect 1642 2056 1644 2064
rect 1652 2056 1654 2064
rect 1642 2054 1654 2056
rect 1770 2064 1782 2066
rect 1770 2056 1772 2064
rect 1780 2056 1782 2064
rect 1576 2006 1578 2014
rect 1586 2006 1590 2014
rect 1598 2006 1602 2014
rect 1610 2006 1614 2014
rect 1622 2006 1624 2014
rect 1482 1944 1494 1946
rect 1482 1936 1484 1944
rect 1492 1936 1494 1944
rect 1482 1884 1494 1936
rect 1482 1876 1484 1884
rect 1492 1876 1494 1884
rect 1482 1874 1494 1876
rect 1546 1824 1558 1826
rect 1546 1816 1548 1824
rect 1556 1816 1558 1824
rect 1514 1764 1526 1766
rect 1514 1756 1516 1764
rect 1524 1756 1526 1764
rect 1450 1496 1452 1504
rect 1460 1496 1462 1504
rect 1450 1494 1462 1496
rect 1482 1524 1494 1526
rect 1482 1516 1484 1524
rect 1492 1516 1494 1524
rect 1418 1456 1420 1464
rect 1428 1456 1430 1464
rect 1418 1454 1430 1456
rect 1386 1356 1388 1364
rect 1396 1356 1398 1364
rect 1386 1354 1398 1356
rect 1418 1364 1430 1366
rect 1418 1356 1420 1364
rect 1428 1356 1430 1364
rect 1354 1304 1366 1306
rect 1354 1296 1356 1304
rect 1364 1296 1366 1304
rect 1354 1044 1366 1296
rect 1354 1036 1356 1044
rect 1364 1036 1366 1044
rect 1354 1034 1366 1036
rect 1386 964 1398 966
rect 1386 956 1388 964
rect 1396 956 1398 964
rect 1386 884 1398 956
rect 1386 876 1388 884
rect 1396 876 1398 884
rect 1386 874 1398 876
rect 1418 846 1430 1356
rect 1482 1364 1494 1516
rect 1514 1424 1526 1756
rect 1546 1684 1558 1816
rect 1546 1676 1548 1684
rect 1556 1676 1558 1684
rect 1546 1674 1558 1676
rect 1576 1614 1624 2006
rect 1674 2004 1686 2006
rect 1674 1996 1676 2004
rect 1684 1996 1686 2004
rect 1674 1864 1686 1996
rect 1706 2004 1718 2006
rect 1706 1996 1708 2004
rect 1716 1996 1718 2004
rect 1706 1884 1718 1996
rect 1706 1876 1708 1884
rect 1716 1876 1718 1884
rect 1706 1874 1718 1876
rect 1738 1924 1750 1926
rect 1738 1916 1740 1924
rect 1748 1916 1750 1924
rect 1674 1856 1676 1864
rect 1684 1856 1686 1864
rect 1674 1854 1686 1856
rect 1642 1824 1654 1826
rect 1642 1816 1644 1824
rect 1652 1816 1654 1824
rect 1642 1806 1654 1816
rect 1738 1824 1750 1916
rect 1738 1816 1740 1824
rect 1748 1816 1750 1824
rect 1738 1814 1750 1816
rect 1642 1794 1686 1806
rect 1576 1606 1578 1614
rect 1586 1606 1590 1614
rect 1598 1606 1602 1614
rect 1610 1606 1614 1614
rect 1622 1606 1624 1614
rect 1514 1416 1516 1424
rect 1524 1416 1526 1424
rect 1514 1414 1526 1416
rect 1546 1544 1558 1546
rect 1546 1536 1548 1544
rect 1556 1536 1558 1544
rect 1482 1356 1484 1364
rect 1492 1356 1494 1364
rect 1482 1354 1494 1356
rect 1546 1364 1558 1536
rect 1546 1356 1548 1364
rect 1556 1356 1558 1364
rect 1546 1354 1558 1356
rect 1482 1324 1494 1326
rect 1482 1316 1484 1324
rect 1492 1316 1494 1324
rect 1482 1264 1494 1316
rect 1482 1256 1484 1264
rect 1492 1256 1494 1264
rect 1482 1254 1494 1256
rect 1514 1224 1526 1226
rect 1514 1216 1516 1224
rect 1524 1216 1526 1224
rect 1450 1124 1462 1126
rect 1450 1116 1452 1124
rect 1460 1116 1462 1124
rect 1450 984 1462 1116
rect 1450 976 1452 984
rect 1460 976 1462 984
rect 1450 974 1462 976
rect 1482 1084 1494 1086
rect 1482 1076 1484 1084
rect 1492 1076 1494 1084
rect 1482 964 1494 1076
rect 1482 956 1484 964
rect 1492 956 1494 964
rect 1482 954 1494 956
rect 1514 1004 1526 1216
rect 1576 1214 1624 1606
rect 1642 1544 1654 1546
rect 1642 1536 1644 1544
rect 1652 1536 1654 1544
rect 1642 1504 1654 1536
rect 1642 1496 1644 1504
rect 1652 1496 1654 1504
rect 1642 1494 1654 1496
rect 1674 1404 1686 1794
rect 1674 1396 1676 1404
rect 1684 1396 1686 1404
rect 1674 1394 1686 1396
rect 1706 1724 1718 1726
rect 1706 1716 1708 1724
rect 1716 1716 1718 1724
rect 1706 1304 1718 1716
rect 1738 1544 1750 1546
rect 1738 1536 1740 1544
rect 1748 1536 1750 1544
rect 1738 1324 1750 1536
rect 1770 1444 1782 2056
rect 1770 1436 1772 1444
rect 1780 1436 1782 1444
rect 1770 1434 1782 1436
rect 1738 1316 1740 1324
rect 1748 1316 1750 1324
rect 1738 1314 1750 1316
rect 1706 1296 1708 1304
rect 1716 1296 1718 1304
rect 1706 1294 1718 1296
rect 1576 1206 1578 1214
rect 1586 1206 1590 1214
rect 1598 1206 1602 1214
rect 1610 1206 1614 1214
rect 1622 1206 1624 1214
rect 1514 996 1516 1004
rect 1524 996 1526 1004
rect 1514 846 1526 996
rect 1546 1004 1558 1006
rect 1546 996 1548 1004
rect 1556 996 1558 1004
rect 1546 904 1558 996
rect 1546 896 1548 904
rect 1556 896 1558 904
rect 1546 894 1558 896
rect 1322 836 1324 844
rect 1332 836 1334 844
rect 1322 834 1334 836
rect 1386 834 1430 846
rect 1482 834 1526 846
rect 1386 804 1398 834
rect 1386 796 1388 804
rect 1396 796 1398 804
rect 1386 794 1398 796
rect 1418 804 1430 806
rect 1418 796 1420 804
rect 1428 796 1430 804
rect 1418 766 1430 796
rect 1354 754 1430 766
rect 1450 764 1462 766
rect 1450 756 1452 764
rect 1460 756 1462 764
rect 1322 744 1334 746
rect 1322 736 1324 744
rect 1332 736 1334 744
rect 1258 704 1270 706
rect 1258 696 1260 704
rect 1268 696 1270 704
rect 1258 664 1270 696
rect 1258 656 1260 664
rect 1268 656 1270 664
rect 1258 654 1270 656
rect 1322 544 1334 736
rect 1322 536 1324 544
rect 1332 536 1334 544
rect 1322 504 1334 536
rect 1322 496 1324 504
rect 1332 496 1334 504
rect 1322 494 1334 496
rect 1322 404 1334 406
rect 1322 396 1324 404
rect 1332 396 1334 404
rect 1258 314 1302 326
rect 1258 284 1270 314
rect 1290 308 1302 314
rect 1290 300 1292 308
rect 1300 300 1302 308
rect 1290 294 1302 300
rect 1322 324 1334 396
rect 1322 316 1324 324
rect 1332 316 1334 324
rect 1258 276 1260 284
rect 1268 276 1270 284
rect 1258 274 1270 276
rect 1290 280 1302 286
rect 1226 256 1228 264
rect 1236 256 1238 264
rect 1226 254 1238 256
rect 1290 272 1292 280
rect 1300 272 1302 280
rect 1162 116 1164 124
rect 1172 116 1174 124
rect 1162 114 1174 116
rect 1258 164 1270 166
rect 1258 156 1260 164
rect 1268 156 1270 164
rect 1258 124 1270 156
rect 1258 116 1260 124
rect 1268 116 1270 124
rect 1258 114 1270 116
rect 938 96 940 104
rect 948 96 950 104
rect 938 94 950 96
rect 1290 104 1302 272
rect 1322 244 1334 316
rect 1354 284 1366 754
rect 1450 604 1462 756
rect 1450 596 1452 604
rect 1460 596 1462 604
rect 1450 594 1462 596
rect 1482 504 1494 834
rect 1576 814 1624 1206
rect 1674 1224 1686 1226
rect 1674 1216 1676 1224
rect 1684 1216 1686 1224
rect 1674 1144 1686 1216
rect 1802 1204 1814 2076
rect 1834 1864 1846 2176
rect 1930 2184 1942 2434
rect 1962 2284 1974 2636
rect 2026 2644 2038 3056
rect 2026 2636 2028 2644
rect 2036 2636 2038 2644
rect 2026 2634 2038 2636
rect 2026 2544 2038 2546
rect 2026 2536 2028 2544
rect 2036 2536 2038 2544
rect 1962 2276 1964 2284
rect 1972 2276 1974 2284
rect 1962 2274 1974 2276
rect 1994 2504 2006 2506
rect 1994 2496 1996 2504
rect 2004 2496 2006 2504
rect 1930 2176 1932 2184
rect 1940 2176 1942 2184
rect 1930 2174 1942 2176
rect 1866 2164 1878 2166
rect 1866 2156 1868 2164
rect 1876 2156 1878 2164
rect 1866 1984 1878 2156
rect 1866 1976 1868 1984
rect 1876 1976 1878 1984
rect 1866 1974 1878 1976
rect 1930 2144 1942 2146
rect 1930 2136 1932 2144
rect 1940 2136 1942 2144
rect 1898 1944 1910 1946
rect 1898 1936 1900 1944
rect 1908 1936 1910 1944
rect 1834 1856 1836 1864
rect 1844 1856 1846 1864
rect 1834 1854 1846 1856
rect 1866 1904 1878 1906
rect 1866 1896 1868 1904
rect 1876 1896 1878 1904
rect 1834 1824 1846 1826
rect 1834 1816 1836 1824
rect 1844 1816 1846 1824
rect 1834 1724 1846 1816
rect 1834 1716 1836 1724
rect 1844 1716 1846 1724
rect 1834 1714 1846 1716
rect 1866 1704 1878 1896
rect 1898 1864 1910 1936
rect 1930 1944 1942 2136
rect 1994 2104 2006 2496
rect 2026 2204 2038 2536
rect 2058 2504 2070 3136
rect 2090 2884 2102 3176
rect 2122 3104 2134 3236
rect 2122 3096 2124 3104
rect 2132 3096 2134 3104
rect 2122 3094 2134 3096
rect 2154 3104 2166 3106
rect 2154 3096 2156 3104
rect 2164 3096 2166 3104
rect 2154 3044 2166 3096
rect 2154 3036 2156 3044
rect 2164 3036 2166 3044
rect 2154 3034 2166 3036
rect 2186 3024 2198 3496
rect 2218 3484 2230 3486
rect 2218 3476 2220 3484
rect 2228 3476 2230 3484
rect 2218 3204 2230 3476
rect 2250 3484 2262 3676
rect 2250 3476 2252 3484
rect 2260 3476 2262 3484
rect 2250 3474 2262 3476
rect 2218 3196 2220 3204
rect 2228 3196 2230 3204
rect 2218 3194 2230 3196
rect 2250 3344 2262 3346
rect 2250 3336 2252 3344
rect 2260 3336 2262 3344
rect 2186 3016 2188 3024
rect 2196 3016 2198 3024
rect 2186 3014 2198 3016
rect 2090 2876 2092 2884
rect 2100 2876 2102 2884
rect 2090 2874 2102 2876
rect 2154 3004 2166 3006
rect 2154 2996 2156 3004
rect 2164 2996 2166 3004
rect 2154 2804 2166 2996
rect 2154 2796 2156 2804
rect 2164 2796 2166 2804
rect 2154 2764 2166 2796
rect 2154 2756 2156 2764
rect 2164 2756 2166 2764
rect 2154 2754 2166 2756
rect 2186 2944 2198 2946
rect 2186 2936 2188 2944
rect 2196 2936 2198 2944
rect 2122 2724 2134 2726
rect 2122 2716 2124 2724
rect 2132 2716 2134 2724
rect 2122 2624 2134 2716
rect 2186 2724 2198 2936
rect 2186 2716 2188 2724
rect 2196 2716 2198 2724
rect 2186 2714 2198 2716
rect 2218 2944 2230 2946
rect 2218 2936 2220 2944
rect 2228 2936 2230 2944
rect 2218 2704 2230 2936
rect 2218 2696 2220 2704
rect 2228 2696 2230 2704
rect 2218 2694 2230 2696
rect 2250 2864 2262 3336
rect 2282 3224 2294 3696
rect 2314 3544 2326 3716
rect 2346 3664 2358 4176
rect 2378 4184 2390 4436
rect 2410 4224 2422 4616
rect 2730 4624 2742 4626
rect 2730 4616 2732 4624
rect 2740 4616 2742 4624
rect 2538 4564 2550 4566
rect 2538 4556 2540 4564
rect 2548 4556 2550 4564
rect 2410 4216 2412 4224
rect 2420 4216 2422 4224
rect 2410 4214 2422 4216
rect 2442 4324 2454 4326
rect 2442 4316 2444 4324
rect 2452 4316 2454 4324
rect 2378 4176 2380 4184
rect 2388 4176 2390 4184
rect 2378 4174 2390 4176
rect 2410 4124 2422 4126
rect 2410 4116 2412 4124
rect 2420 4116 2422 4124
rect 2378 4104 2390 4106
rect 2378 4096 2380 4104
rect 2388 4096 2390 4104
rect 2378 4044 2390 4096
rect 2378 4036 2380 4044
rect 2388 4036 2390 4044
rect 2378 3904 2390 4036
rect 2378 3896 2380 3904
rect 2388 3896 2390 3904
rect 2378 3894 2390 3896
rect 2410 4084 2422 4116
rect 2442 4124 2454 4316
rect 2442 4116 2444 4124
rect 2452 4116 2454 4124
rect 2442 4114 2454 4116
rect 2506 4244 2518 4246
rect 2506 4236 2508 4244
rect 2516 4236 2518 4244
rect 2506 4104 2518 4236
rect 2506 4096 2508 4104
rect 2516 4096 2518 4104
rect 2506 4094 2518 4096
rect 2410 4076 2412 4084
rect 2420 4076 2422 4084
rect 2346 3656 2348 3664
rect 2356 3656 2358 3664
rect 2346 3654 2358 3656
rect 2378 3684 2390 3686
rect 2378 3676 2380 3684
rect 2388 3676 2390 3684
rect 2314 3536 2316 3544
rect 2324 3536 2326 3544
rect 2314 3534 2326 3536
rect 2346 3524 2358 3526
rect 2346 3516 2348 3524
rect 2356 3516 2358 3524
rect 2314 3424 2326 3426
rect 2314 3416 2316 3424
rect 2324 3416 2326 3424
rect 2314 3364 2326 3416
rect 2314 3356 2316 3364
rect 2324 3356 2326 3364
rect 2314 3354 2326 3356
rect 2346 3264 2358 3516
rect 2378 3344 2390 3676
rect 2410 3584 2422 4076
rect 2442 3984 2454 3986
rect 2442 3976 2444 3984
rect 2452 3976 2454 3984
rect 2442 3944 2454 3976
rect 2442 3936 2444 3944
rect 2452 3936 2454 3944
rect 2442 3934 2454 3936
rect 2474 3964 2486 3966
rect 2474 3956 2476 3964
rect 2484 3956 2486 3964
rect 2442 3744 2454 3746
rect 2442 3736 2444 3744
rect 2452 3736 2454 3744
rect 2442 3684 2454 3736
rect 2442 3676 2444 3684
rect 2452 3676 2454 3684
rect 2442 3674 2454 3676
rect 2410 3576 2412 3584
rect 2420 3576 2422 3584
rect 2410 3574 2422 3576
rect 2442 3564 2454 3566
rect 2442 3556 2444 3564
rect 2452 3556 2454 3564
rect 2410 3504 2422 3506
rect 2410 3496 2412 3504
rect 2420 3496 2422 3504
rect 2410 3404 2422 3496
rect 2410 3396 2412 3404
rect 2420 3396 2422 3404
rect 2410 3394 2422 3396
rect 2378 3336 2380 3344
rect 2388 3336 2390 3344
rect 2378 3334 2390 3336
rect 2410 3344 2422 3346
rect 2410 3336 2412 3344
rect 2420 3336 2422 3344
rect 2346 3256 2348 3264
rect 2356 3256 2358 3264
rect 2346 3254 2358 3256
rect 2282 3216 2284 3224
rect 2292 3216 2294 3224
rect 2282 3214 2294 3216
rect 2378 3084 2390 3086
rect 2378 3076 2380 3084
rect 2388 3076 2390 3084
rect 2346 3064 2358 3066
rect 2346 3056 2348 3064
rect 2356 3056 2358 3064
rect 2282 3024 2294 3026
rect 2282 3016 2284 3024
rect 2292 3016 2294 3024
rect 2282 2904 2294 3016
rect 2282 2896 2284 2904
rect 2292 2896 2294 2904
rect 2282 2894 2294 2896
rect 2346 2884 2358 3056
rect 2346 2876 2348 2884
rect 2356 2876 2358 2884
rect 2346 2874 2358 2876
rect 2250 2856 2252 2864
rect 2260 2856 2262 2864
rect 2122 2616 2124 2624
rect 2132 2616 2134 2624
rect 2122 2614 2134 2616
rect 2186 2684 2198 2686
rect 2186 2676 2188 2684
rect 2196 2676 2198 2684
rect 2186 2544 2198 2676
rect 2250 2664 2262 2856
rect 2250 2656 2252 2664
rect 2260 2656 2262 2664
rect 2250 2654 2262 2656
rect 2346 2764 2358 2766
rect 2346 2756 2348 2764
rect 2356 2756 2358 2764
rect 2346 2664 2358 2756
rect 2346 2656 2348 2664
rect 2356 2656 2358 2664
rect 2346 2654 2358 2656
rect 2378 2764 2390 3076
rect 2378 2756 2380 2764
rect 2388 2756 2390 2764
rect 2250 2624 2262 2626
rect 2250 2616 2252 2624
rect 2260 2616 2262 2624
rect 2186 2536 2188 2544
rect 2196 2536 2198 2544
rect 2186 2534 2198 2536
rect 2218 2604 2230 2606
rect 2218 2596 2220 2604
rect 2228 2596 2230 2604
rect 2058 2496 2060 2504
rect 2068 2496 2070 2504
rect 2058 2494 2070 2496
rect 2090 2524 2102 2526
rect 2090 2516 2092 2524
rect 2100 2516 2102 2524
rect 2090 2484 2102 2516
rect 2090 2476 2092 2484
rect 2100 2476 2102 2484
rect 2090 2474 2102 2476
rect 2154 2504 2166 2506
rect 2154 2496 2156 2504
rect 2164 2496 2166 2504
rect 2058 2424 2070 2426
rect 2058 2416 2060 2424
rect 2068 2416 2070 2424
rect 2058 2364 2070 2416
rect 2058 2356 2060 2364
rect 2068 2356 2070 2364
rect 2058 2354 2070 2356
rect 2090 2404 2102 2406
rect 2090 2396 2092 2404
rect 2100 2396 2102 2404
rect 2090 2264 2102 2396
rect 2090 2256 2092 2264
rect 2100 2256 2102 2264
rect 2090 2254 2102 2256
rect 2122 2344 2134 2346
rect 2122 2336 2124 2344
rect 2132 2336 2134 2344
rect 2026 2196 2028 2204
rect 2036 2196 2038 2204
rect 2026 2194 2038 2196
rect 2122 2164 2134 2336
rect 2122 2156 2124 2164
rect 2132 2156 2134 2164
rect 2122 2154 2134 2156
rect 2154 2144 2166 2496
rect 2218 2364 2230 2596
rect 2250 2404 2262 2616
rect 2314 2544 2326 2546
rect 2314 2536 2316 2544
rect 2324 2536 2326 2544
rect 2250 2396 2252 2404
rect 2260 2396 2262 2404
rect 2250 2394 2262 2396
rect 2282 2404 2294 2406
rect 2282 2396 2284 2404
rect 2292 2396 2294 2404
rect 2218 2356 2220 2364
rect 2228 2356 2230 2364
rect 2218 2354 2230 2356
rect 2218 2324 2230 2326
rect 2218 2316 2220 2324
rect 2228 2316 2230 2324
rect 2154 2136 2156 2144
rect 2164 2136 2166 2144
rect 2154 2134 2166 2136
rect 2186 2264 2198 2266
rect 2186 2256 2188 2264
rect 2196 2256 2198 2264
rect 1994 2096 1996 2104
rect 2004 2096 2006 2104
rect 1994 2094 2006 2096
rect 2058 2104 2070 2106
rect 2058 2096 2060 2104
rect 2068 2096 2070 2104
rect 2058 2086 2070 2096
rect 1978 2084 2070 2086
rect 1978 2076 1980 2084
rect 1988 2076 2070 2084
rect 1978 2074 2070 2076
rect 2154 2104 2166 2106
rect 2154 2096 2156 2104
rect 2164 2096 2166 2104
rect 1930 1936 1932 1944
rect 1940 1936 1942 1944
rect 1930 1934 1942 1936
rect 1962 2004 1974 2006
rect 1962 1996 1964 2004
rect 1972 1996 1974 2004
rect 1898 1856 1900 1864
rect 1908 1856 1910 1864
rect 1898 1854 1910 1856
rect 1930 1904 1942 1906
rect 1930 1896 1932 1904
rect 1940 1896 1942 1904
rect 1866 1696 1868 1704
rect 1876 1696 1878 1704
rect 1866 1694 1878 1696
rect 1898 1724 1910 1726
rect 1898 1716 1900 1724
rect 1908 1716 1910 1724
rect 1866 1584 1878 1586
rect 1866 1576 1868 1584
rect 1876 1576 1878 1584
rect 1834 1544 1846 1546
rect 1834 1536 1836 1544
rect 1844 1536 1846 1544
rect 1834 1404 1846 1536
rect 1866 1484 1878 1576
rect 1866 1476 1868 1484
rect 1876 1476 1878 1484
rect 1866 1474 1878 1476
rect 1834 1396 1836 1404
rect 1844 1396 1846 1404
rect 1834 1394 1846 1396
rect 1802 1196 1804 1204
rect 1812 1196 1814 1204
rect 1802 1194 1814 1196
rect 1834 1364 1846 1366
rect 1834 1356 1836 1364
rect 1844 1356 1846 1364
rect 1674 1136 1676 1144
rect 1684 1136 1686 1144
rect 1674 1134 1686 1136
rect 1706 1124 1718 1126
rect 1706 1116 1708 1124
rect 1716 1116 1718 1124
rect 1642 1044 1654 1046
rect 1642 1036 1644 1044
rect 1652 1036 1654 1044
rect 1642 904 1654 1036
rect 1706 1044 1718 1116
rect 1834 1124 1846 1356
rect 1834 1116 1836 1124
rect 1844 1116 1846 1124
rect 1834 1114 1846 1116
rect 1706 1036 1708 1044
rect 1716 1036 1718 1044
rect 1706 1034 1718 1036
rect 1802 1084 1814 1086
rect 1802 1076 1804 1084
rect 1812 1076 1814 1084
rect 1642 896 1644 904
rect 1652 896 1654 904
rect 1642 894 1654 896
rect 1770 924 1782 926
rect 1770 916 1772 924
rect 1780 916 1782 924
rect 1576 806 1578 814
rect 1586 806 1590 814
rect 1598 806 1602 814
rect 1610 806 1614 814
rect 1622 806 1624 814
rect 1514 784 1526 786
rect 1514 776 1516 784
rect 1524 776 1526 784
rect 1514 584 1526 776
rect 1514 576 1516 584
rect 1524 576 1526 584
rect 1514 574 1526 576
rect 1482 496 1484 504
rect 1492 496 1494 504
rect 1482 494 1494 496
rect 1576 414 1624 806
rect 1674 804 1686 806
rect 1674 796 1676 804
rect 1684 796 1686 804
rect 1674 544 1686 796
rect 1738 804 1750 806
rect 1738 796 1740 804
rect 1748 796 1750 804
rect 1738 644 1750 796
rect 1770 664 1782 916
rect 1802 924 1814 1076
rect 1866 1084 1878 1086
rect 1866 1076 1868 1084
rect 1876 1076 1878 1084
rect 1802 916 1804 924
rect 1812 916 1814 924
rect 1802 914 1814 916
rect 1834 1044 1846 1046
rect 1834 1036 1836 1044
rect 1844 1036 1846 1044
rect 1834 764 1846 1036
rect 1866 964 1878 1076
rect 1866 956 1868 964
rect 1876 956 1878 964
rect 1866 954 1878 956
rect 1834 756 1836 764
rect 1844 756 1846 764
rect 1834 754 1846 756
rect 1866 904 1878 906
rect 1866 896 1868 904
rect 1876 896 1878 904
rect 1866 764 1878 896
rect 1866 756 1868 764
rect 1876 756 1878 764
rect 1866 754 1878 756
rect 1898 784 1910 1716
rect 1930 1606 1942 1896
rect 1962 1724 1974 1996
rect 1994 1984 2006 1986
rect 1994 1976 1996 1984
rect 2004 1976 2006 1984
rect 1994 1864 2006 1976
rect 2090 1984 2102 1986
rect 2090 1976 2092 1984
rect 2100 1976 2102 1984
rect 1994 1856 1996 1864
rect 2004 1856 2006 1864
rect 1994 1854 2006 1856
rect 2026 1904 2038 1906
rect 2026 1896 2028 1904
rect 2036 1896 2038 1904
rect 1962 1716 1964 1724
rect 1972 1716 1974 1724
rect 1962 1714 1974 1716
rect 1994 1764 2006 1766
rect 1994 1756 1996 1764
rect 2004 1756 2006 1764
rect 1994 1684 2006 1756
rect 1994 1676 1996 1684
rect 2004 1676 2006 1684
rect 1994 1674 2006 1676
rect 1914 1604 1942 1606
rect 1914 1596 1916 1604
rect 1924 1596 1942 1604
rect 1914 1594 1942 1596
rect 1994 1644 2006 1646
rect 1994 1636 1996 1644
rect 2004 1636 2006 1644
rect 1962 1584 1974 1586
rect 1962 1576 1964 1584
rect 1972 1576 1974 1584
rect 1930 1524 1942 1526
rect 1930 1516 1932 1524
rect 1940 1516 1942 1524
rect 1930 1084 1942 1516
rect 1962 1324 1974 1576
rect 1962 1316 1964 1324
rect 1972 1316 1974 1324
rect 1962 1314 1974 1316
rect 1962 1284 1974 1286
rect 1962 1276 1964 1284
rect 1972 1276 1974 1284
rect 1962 1104 1974 1276
rect 1962 1096 1964 1104
rect 1972 1096 1974 1104
rect 1962 1094 1974 1096
rect 1930 1076 1932 1084
rect 1940 1076 1942 1084
rect 1930 1074 1942 1076
rect 1962 1044 1974 1046
rect 1962 1036 1964 1044
rect 1972 1036 1974 1044
rect 1962 1004 1974 1036
rect 1962 996 1964 1004
rect 1972 996 1974 1004
rect 1962 994 1974 996
rect 1994 964 2006 1636
rect 2026 1304 2038 1896
rect 2058 1904 2070 1906
rect 2058 1896 2060 1904
rect 2068 1896 2070 1904
rect 2058 1744 2070 1896
rect 2090 1884 2102 1976
rect 2090 1876 2092 1884
rect 2100 1876 2102 1884
rect 2090 1874 2102 1876
rect 2122 1944 2134 1946
rect 2122 1936 2124 1944
rect 2132 1936 2134 1944
rect 2058 1736 2060 1744
rect 2068 1736 2070 1744
rect 2058 1734 2070 1736
rect 2090 1844 2102 1846
rect 2090 1836 2092 1844
rect 2100 1836 2102 1844
rect 2058 1664 2070 1666
rect 2058 1656 2060 1664
rect 2068 1656 2070 1664
rect 2058 1504 2070 1656
rect 2090 1524 2102 1836
rect 2122 1804 2134 1936
rect 2154 1924 2166 2096
rect 2154 1916 2156 1924
rect 2164 1916 2166 1924
rect 2154 1914 2166 1916
rect 2186 1904 2198 2256
rect 2218 2104 2230 2316
rect 2250 2304 2262 2306
rect 2250 2296 2252 2304
rect 2260 2296 2262 2304
rect 2250 2184 2262 2296
rect 2250 2176 2252 2184
rect 2260 2176 2262 2184
rect 2250 2174 2262 2176
rect 2282 2184 2294 2396
rect 2314 2404 2326 2536
rect 2314 2396 2316 2404
rect 2324 2396 2326 2404
rect 2314 2394 2326 2396
rect 2378 2384 2390 2756
rect 2410 2544 2422 3336
rect 2442 3164 2454 3556
rect 2474 3504 2486 3956
rect 2538 3924 2550 4556
rect 2698 4524 2710 4526
rect 2698 4516 2700 4524
rect 2708 4516 2710 4524
rect 2570 4444 2582 4446
rect 2570 4436 2572 4444
rect 2580 4436 2582 4444
rect 2570 4084 2582 4436
rect 2570 4076 2572 4084
rect 2580 4076 2582 4084
rect 2570 4074 2582 4076
rect 2634 4164 2646 4166
rect 2634 4156 2636 4164
rect 2644 4156 2646 4164
rect 2538 3916 2540 3924
rect 2548 3916 2550 3924
rect 2538 3914 2550 3916
rect 2570 4044 2582 4046
rect 2570 4036 2572 4044
rect 2580 4036 2582 4044
rect 2570 3884 2582 4036
rect 2634 4024 2646 4156
rect 2634 4016 2636 4024
rect 2644 4016 2646 4024
rect 2634 4014 2646 4016
rect 2666 4124 2678 4126
rect 2666 4116 2668 4124
rect 2676 4116 2678 4124
rect 2570 3876 2572 3884
rect 2580 3876 2582 3884
rect 2570 3874 2582 3876
rect 2602 3984 2614 3986
rect 2602 3976 2604 3984
rect 2612 3976 2614 3984
rect 2506 3784 2518 3786
rect 2506 3776 2508 3784
rect 2516 3776 2518 3784
rect 2506 3684 2518 3776
rect 2506 3676 2508 3684
rect 2516 3676 2518 3684
rect 2506 3674 2518 3676
rect 2538 3784 2550 3786
rect 2538 3776 2540 3784
rect 2548 3776 2550 3784
rect 2474 3496 2476 3504
rect 2484 3496 2486 3504
rect 2474 3494 2486 3496
rect 2506 3604 2518 3606
rect 2506 3596 2508 3604
rect 2516 3596 2518 3604
rect 2442 3156 2444 3164
rect 2452 3156 2454 3164
rect 2442 3154 2454 3156
rect 2474 3404 2486 3406
rect 2474 3396 2476 3404
rect 2484 3396 2486 3404
rect 2442 3124 2454 3126
rect 2442 3116 2444 3124
rect 2452 3116 2454 3124
rect 2442 3064 2454 3116
rect 2474 3104 2486 3396
rect 2506 3224 2518 3596
rect 2538 3564 2550 3776
rect 2602 3704 2614 3976
rect 2602 3696 2604 3704
rect 2612 3696 2614 3704
rect 2602 3694 2614 3696
rect 2634 3944 2646 3946
rect 2634 3936 2636 3944
rect 2644 3936 2646 3944
rect 2602 3644 2614 3646
rect 2602 3636 2604 3644
rect 2612 3636 2614 3644
rect 2538 3556 2540 3564
rect 2548 3556 2550 3564
rect 2538 3554 2550 3556
rect 2570 3604 2582 3606
rect 2570 3596 2572 3604
rect 2580 3596 2582 3604
rect 2570 3364 2582 3596
rect 2570 3356 2572 3364
rect 2580 3356 2582 3364
rect 2506 3216 2508 3224
rect 2516 3216 2518 3224
rect 2506 3214 2518 3216
rect 2538 3324 2550 3326
rect 2538 3316 2540 3324
rect 2548 3316 2550 3324
rect 2474 3096 2476 3104
rect 2484 3096 2486 3104
rect 2474 3094 2486 3096
rect 2506 3164 2518 3166
rect 2506 3156 2508 3164
rect 2516 3156 2518 3164
rect 2506 3084 2518 3156
rect 2506 3076 2508 3084
rect 2516 3076 2518 3084
rect 2506 3074 2518 3076
rect 2442 3056 2444 3064
rect 2452 3056 2454 3064
rect 2442 3054 2454 3056
rect 2538 3044 2550 3316
rect 2538 3036 2540 3044
rect 2548 3036 2550 3044
rect 2538 3034 2550 3036
rect 2570 3204 2582 3356
rect 2570 3196 2572 3204
rect 2580 3196 2582 3204
rect 2506 3024 2518 3026
rect 2506 3016 2508 3024
rect 2516 3016 2518 3024
rect 2474 2964 2486 2966
rect 2474 2956 2476 2964
rect 2484 2956 2486 2964
rect 2442 2944 2454 2946
rect 2442 2936 2444 2944
rect 2452 2936 2454 2944
rect 2442 2824 2454 2936
rect 2442 2816 2444 2824
rect 2452 2816 2454 2824
rect 2442 2814 2454 2816
rect 2410 2536 2412 2544
rect 2420 2536 2422 2544
rect 2410 2534 2422 2536
rect 2442 2684 2454 2686
rect 2442 2676 2444 2684
rect 2452 2676 2454 2684
rect 2394 2484 2422 2486
rect 2394 2476 2396 2484
rect 2404 2476 2422 2484
rect 2394 2474 2422 2476
rect 2378 2376 2380 2384
rect 2388 2376 2390 2384
rect 2378 2374 2390 2376
rect 2378 2304 2390 2306
rect 2378 2296 2380 2304
rect 2388 2296 2390 2304
rect 2282 2176 2284 2184
rect 2292 2176 2294 2184
rect 2282 2174 2294 2176
rect 2314 2264 2326 2266
rect 2314 2256 2316 2264
rect 2324 2256 2326 2264
rect 2218 2096 2220 2104
rect 2228 2096 2230 2104
rect 2218 2094 2230 2096
rect 2250 1984 2262 1986
rect 2250 1976 2252 1984
rect 2260 1976 2262 1984
rect 2186 1896 2188 1904
rect 2196 1896 2198 1904
rect 2186 1894 2198 1896
rect 2218 1944 2230 1946
rect 2218 1936 2220 1944
rect 2228 1936 2230 1944
rect 2154 1884 2166 1886
rect 2154 1876 2156 1884
rect 2164 1876 2166 1884
rect 2154 1824 2166 1876
rect 2154 1816 2156 1824
rect 2164 1816 2166 1824
rect 2154 1814 2166 1816
rect 2122 1796 2124 1804
rect 2132 1796 2134 1804
rect 2122 1794 2134 1796
rect 2186 1804 2198 1806
rect 2186 1796 2188 1804
rect 2196 1796 2198 1804
rect 2154 1744 2166 1746
rect 2154 1736 2156 1744
rect 2164 1736 2166 1744
rect 2154 1704 2166 1736
rect 2154 1696 2156 1704
rect 2164 1696 2166 1704
rect 2154 1694 2166 1696
rect 2090 1516 2092 1524
rect 2100 1516 2102 1524
rect 2090 1514 2102 1516
rect 2122 1544 2134 1546
rect 2122 1536 2124 1544
rect 2132 1536 2134 1544
rect 2058 1496 2060 1504
rect 2068 1496 2070 1504
rect 2058 1494 2070 1496
rect 2090 1484 2102 1486
rect 2090 1476 2092 1484
rect 2100 1476 2102 1484
rect 2026 1296 2028 1304
rect 2036 1296 2038 1304
rect 2026 1294 2038 1296
rect 2058 1444 2070 1446
rect 2058 1436 2060 1444
rect 2068 1436 2070 1444
rect 2058 1304 2070 1436
rect 2090 1324 2102 1476
rect 2090 1316 2092 1324
rect 2100 1316 2102 1324
rect 2090 1314 2102 1316
rect 2058 1296 2060 1304
rect 2068 1296 2070 1304
rect 1994 956 1996 964
rect 2004 956 2006 964
rect 1994 954 2006 956
rect 2058 924 2070 1296
rect 2122 1284 2134 1536
rect 2122 1276 2124 1284
rect 2132 1276 2134 1284
rect 2122 1274 2134 1276
rect 2154 1464 2166 1466
rect 2154 1456 2156 1464
rect 2164 1456 2166 1464
rect 2090 1264 2102 1266
rect 2090 1256 2092 1264
rect 2100 1256 2102 1264
rect 2090 984 2102 1256
rect 2154 1184 2166 1456
rect 2186 1464 2198 1796
rect 2218 1684 2230 1936
rect 2250 1864 2262 1976
rect 2314 1886 2326 2256
rect 2346 2204 2358 2206
rect 2346 2196 2348 2204
rect 2356 2196 2358 2204
rect 2346 2164 2358 2196
rect 2346 2156 2348 2164
rect 2356 2156 2358 2164
rect 2346 2154 2358 2156
rect 2314 1884 2342 1886
rect 2314 1876 2332 1884
rect 2340 1876 2342 1884
rect 2314 1874 2342 1876
rect 2250 1856 2252 1864
rect 2260 1856 2262 1864
rect 2250 1854 2262 1856
rect 2378 1864 2390 2296
rect 2410 2206 2422 2474
rect 2394 2204 2422 2206
rect 2394 2196 2396 2204
rect 2404 2196 2422 2204
rect 2394 2194 2422 2196
rect 2378 1856 2380 1864
rect 2388 1856 2390 1864
rect 2378 1854 2390 1856
rect 2410 1924 2422 1926
rect 2410 1916 2412 1924
rect 2420 1916 2422 1924
rect 2282 1844 2294 1846
rect 2282 1836 2284 1844
rect 2292 1836 2294 1844
rect 2218 1676 2220 1684
rect 2228 1676 2230 1684
rect 2218 1674 2230 1676
rect 2250 1784 2262 1786
rect 2250 1776 2252 1784
rect 2260 1776 2262 1784
rect 2186 1456 2188 1464
rect 2196 1456 2198 1464
rect 2186 1454 2198 1456
rect 2250 1484 2262 1776
rect 2282 1784 2294 1836
rect 2282 1776 2284 1784
rect 2292 1776 2294 1784
rect 2282 1774 2294 1776
rect 2314 1824 2326 1826
rect 2314 1816 2316 1824
rect 2324 1816 2326 1824
rect 2314 1744 2326 1816
rect 2378 1824 2390 1826
rect 2378 1816 2380 1824
rect 2388 1816 2390 1824
rect 2314 1736 2316 1744
rect 2324 1736 2326 1744
rect 2314 1734 2326 1736
rect 2346 1804 2358 1806
rect 2346 1796 2348 1804
rect 2356 1796 2358 1804
rect 2346 1744 2358 1796
rect 2346 1736 2348 1744
rect 2356 1736 2358 1744
rect 2346 1734 2358 1736
rect 2282 1724 2294 1726
rect 2282 1716 2284 1724
rect 2292 1716 2294 1724
rect 2282 1544 2294 1716
rect 2378 1684 2390 1816
rect 2378 1676 2380 1684
rect 2388 1676 2390 1684
rect 2378 1674 2390 1676
rect 2282 1536 2284 1544
rect 2292 1536 2294 1544
rect 2282 1534 2294 1536
rect 2378 1544 2390 1546
rect 2378 1536 2380 1544
rect 2388 1536 2390 1544
rect 2314 1524 2326 1526
rect 2314 1516 2316 1524
rect 2324 1516 2326 1524
rect 2250 1476 2252 1484
rect 2260 1476 2262 1484
rect 2250 1424 2262 1476
rect 2250 1416 2252 1424
rect 2260 1416 2262 1424
rect 2154 1176 2156 1184
rect 2164 1176 2166 1184
rect 2154 1174 2166 1176
rect 2186 1364 2198 1366
rect 2186 1356 2188 1364
rect 2196 1356 2198 1364
rect 2186 1126 2198 1356
rect 2250 1364 2262 1416
rect 2250 1356 2252 1364
rect 2260 1356 2262 1364
rect 2250 1354 2262 1356
rect 2282 1484 2294 1486
rect 2282 1476 2284 1484
rect 2292 1476 2294 1484
rect 2282 1326 2294 1476
rect 2314 1364 2326 1516
rect 2314 1356 2316 1364
rect 2324 1356 2326 1364
rect 2314 1354 2326 1356
rect 2346 1344 2358 1346
rect 2346 1336 2348 1344
rect 2356 1336 2358 1344
rect 2282 1314 2326 1326
rect 2282 1244 2294 1246
rect 2282 1236 2284 1244
rect 2292 1236 2294 1244
rect 2154 1114 2198 1126
rect 2218 1204 2230 1206
rect 2218 1196 2220 1204
rect 2228 1196 2230 1204
rect 2218 1124 2230 1196
rect 2218 1116 2220 1124
rect 2228 1116 2230 1124
rect 2218 1114 2230 1116
rect 2250 1204 2262 1206
rect 2250 1196 2252 1204
rect 2260 1196 2262 1204
rect 2090 976 2092 984
rect 2100 976 2102 984
rect 2090 974 2102 976
rect 2122 984 2134 986
rect 2122 976 2124 984
rect 2132 976 2134 984
rect 2058 916 2060 924
rect 2068 916 2070 924
rect 2058 914 2070 916
rect 2090 864 2102 866
rect 2090 856 2092 864
rect 2100 856 2102 864
rect 1898 776 1900 784
rect 1908 776 1910 784
rect 1770 656 1772 664
rect 1780 656 1782 664
rect 1770 654 1782 656
rect 1866 724 1878 726
rect 1866 716 1868 724
rect 1876 716 1878 724
rect 1866 646 1878 716
rect 1738 636 1740 644
rect 1748 636 1750 644
rect 1738 634 1750 636
rect 1834 634 1878 646
rect 1834 624 1846 634
rect 1834 616 1836 624
rect 1844 616 1846 624
rect 1834 614 1846 616
rect 1866 624 1878 626
rect 1866 616 1868 624
rect 1876 616 1878 624
rect 1674 536 1676 544
rect 1684 536 1686 544
rect 1674 534 1686 536
rect 1738 584 1750 586
rect 1738 576 1740 584
rect 1748 576 1750 584
rect 1576 406 1578 414
rect 1586 406 1590 414
rect 1598 406 1602 414
rect 1610 406 1614 414
rect 1622 406 1624 414
rect 1482 404 1494 406
rect 1482 396 1484 404
rect 1492 396 1494 404
rect 1482 366 1494 396
rect 1482 354 1526 366
rect 1354 276 1356 284
rect 1364 276 1366 284
rect 1354 274 1366 276
rect 1418 314 1494 326
rect 1418 284 1430 314
rect 1418 276 1420 284
rect 1428 276 1430 284
rect 1418 274 1430 276
rect 1482 284 1494 314
rect 1482 276 1484 284
rect 1492 276 1494 284
rect 1482 274 1494 276
rect 1514 284 1526 354
rect 1514 276 1516 284
rect 1524 276 1526 284
rect 1514 274 1526 276
rect 1322 236 1324 244
rect 1332 236 1334 244
rect 1322 234 1334 236
rect 1530 244 1558 246
rect 1530 236 1532 244
rect 1540 236 1558 244
rect 1530 234 1558 236
rect 1354 204 1366 206
rect 1354 196 1356 204
rect 1364 196 1366 204
rect 1354 164 1366 196
rect 1498 204 1526 206
rect 1498 196 1500 204
rect 1508 196 1526 204
rect 1498 194 1526 196
rect 1354 156 1356 164
rect 1364 156 1366 164
rect 1354 154 1366 156
rect 1514 124 1526 194
rect 1514 116 1516 124
rect 1524 116 1526 124
rect 1514 114 1526 116
rect 1290 96 1292 104
rect 1300 96 1302 104
rect 1290 94 1302 96
rect 1546 64 1558 234
rect 1546 56 1548 64
rect 1556 56 1558 64
rect 1546 54 1558 56
rect 234 36 236 44
rect 244 36 246 44
rect 234 34 246 36
rect 1576 14 1624 406
rect 1674 504 1686 506
rect 1674 496 1676 504
rect 1684 496 1686 504
rect 1674 224 1686 496
rect 1674 216 1676 224
rect 1684 216 1686 224
rect 1674 214 1686 216
rect 1706 284 1718 286
rect 1706 276 1708 284
rect 1716 276 1718 284
rect 1706 166 1718 276
rect 1738 204 1750 576
rect 1802 524 1814 526
rect 1802 516 1804 524
rect 1812 516 1814 524
rect 1802 424 1814 516
rect 1866 446 1878 616
rect 1802 416 1804 424
rect 1812 416 1814 424
rect 1802 414 1814 416
rect 1834 434 1878 446
rect 1770 404 1782 406
rect 1770 396 1772 404
rect 1780 396 1782 404
rect 1770 284 1782 396
rect 1770 276 1772 284
rect 1780 276 1782 284
rect 1770 274 1782 276
rect 1834 206 1846 434
rect 1898 304 1910 776
rect 2058 804 2070 806
rect 2058 796 2060 804
rect 2068 796 2070 804
rect 2026 764 2038 766
rect 2026 756 2028 764
rect 2036 756 2038 764
rect 1962 744 1974 746
rect 1962 736 1964 744
rect 1972 736 1974 744
rect 1930 524 1942 526
rect 1930 516 1932 524
rect 1940 516 1942 524
rect 1930 444 1942 516
rect 1962 524 1974 736
rect 2026 684 2038 756
rect 2026 676 2028 684
rect 2036 676 2038 684
rect 2026 674 2038 676
rect 2058 664 2070 796
rect 2058 656 2060 664
rect 2068 656 2070 664
rect 2058 654 2070 656
rect 1962 516 1964 524
rect 1972 516 1974 524
rect 1962 514 1974 516
rect 1994 624 2006 626
rect 1994 616 1996 624
rect 2004 616 2006 624
rect 1930 436 1932 444
rect 1940 436 1942 444
rect 1930 434 1942 436
rect 1898 296 1900 304
rect 1908 296 1910 304
rect 1898 294 1910 296
rect 1930 364 1942 366
rect 1930 356 1932 364
rect 1940 356 1942 364
rect 1930 304 1942 356
rect 1930 296 1932 304
rect 1940 296 1942 304
rect 1930 294 1942 296
rect 1962 364 1974 366
rect 1962 356 1964 364
rect 1972 356 1974 364
rect 1962 244 1974 356
rect 1994 304 2006 616
rect 2058 624 2070 626
rect 2058 616 2060 624
rect 2068 616 2070 624
rect 1994 296 1996 304
rect 2004 296 2006 304
rect 1994 294 2006 296
rect 2026 544 2038 546
rect 2026 536 2028 544
rect 2036 536 2038 544
rect 1962 236 1964 244
rect 1972 236 1974 244
rect 1962 234 1974 236
rect 1738 196 1740 204
rect 1748 196 1750 204
rect 1738 194 1750 196
rect 1770 204 1782 206
rect 1770 196 1772 204
rect 1780 196 1782 204
rect 1770 166 1782 196
rect 1818 204 1846 206
rect 1818 196 1820 204
rect 1828 196 1846 204
rect 1818 194 1846 196
rect 1898 224 1910 226
rect 1898 216 1900 224
rect 1908 216 1910 224
rect 1706 154 1782 166
rect 1898 124 1910 216
rect 1898 116 1900 124
rect 1908 116 1910 124
rect 1898 114 1910 116
rect 1962 184 1974 186
rect 1962 176 1964 184
rect 1972 176 1974 184
rect 1962 124 1974 176
rect 2026 184 2038 536
rect 2026 176 2028 184
rect 2036 176 2038 184
rect 2026 174 2038 176
rect 2058 144 2070 616
rect 2090 564 2102 856
rect 2122 764 2134 976
rect 2154 804 2166 1114
rect 2154 796 2156 804
rect 2164 796 2166 804
rect 2154 794 2166 796
rect 2186 1084 2198 1086
rect 2186 1076 2188 1084
rect 2196 1076 2198 1084
rect 2186 824 2198 1076
rect 2218 1084 2230 1086
rect 2218 1076 2220 1084
rect 2228 1076 2230 1084
rect 2218 1004 2230 1076
rect 2218 996 2220 1004
rect 2228 996 2230 1004
rect 2218 994 2230 996
rect 2186 816 2188 824
rect 2196 816 2198 824
rect 2122 756 2124 764
rect 2132 756 2134 764
rect 2122 754 2134 756
rect 2186 744 2198 816
rect 2186 736 2188 744
rect 2196 736 2198 744
rect 2186 734 2198 736
rect 2218 964 2230 966
rect 2218 956 2220 964
rect 2228 956 2230 964
rect 2218 744 2230 956
rect 2250 904 2262 1196
rect 2282 1204 2294 1236
rect 2314 1224 2326 1314
rect 2346 1284 2358 1336
rect 2346 1276 2348 1284
rect 2356 1276 2358 1284
rect 2346 1274 2358 1276
rect 2378 1284 2390 1536
rect 2410 1524 2422 1916
rect 2442 1824 2454 2676
rect 2474 2684 2486 2956
rect 2474 2676 2476 2684
rect 2484 2676 2486 2684
rect 2474 2674 2486 2676
rect 2474 2584 2486 2586
rect 2474 2576 2476 2584
rect 2484 2576 2486 2584
rect 2474 2304 2486 2576
rect 2506 2326 2518 3016
rect 2538 3004 2550 3006
rect 2538 2996 2540 3004
rect 2548 2996 2550 3004
rect 2538 2864 2550 2996
rect 2538 2856 2540 2864
rect 2548 2856 2550 2864
rect 2538 2566 2550 2856
rect 2522 2564 2550 2566
rect 2522 2556 2524 2564
rect 2532 2556 2550 2564
rect 2522 2554 2550 2556
rect 2522 2524 2550 2526
rect 2522 2516 2524 2524
rect 2532 2516 2550 2524
rect 2522 2514 2550 2516
rect 2506 2324 2534 2326
rect 2506 2316 2524 2324
rect 2532 2316 2534 2324
rect 2506 2314 2534 2316
rect 2474 2296 2476 2304
rect 2484 2296 2486 2304
rect 2474 2294 2486 2296
rect 2538 2304 2550 2514
rect 2538 2296 2540 2304
rect 2548 2296 2550 2304
rect 2538 2294 2550 2296
rect 2570 2284 2582 3196
rect 2602 3084 2614 3636
rect 2634 3484 2646 3936
rect 2666 3884 2678 4116
rect 2698 3944 2710 4516
rect 2730 4004 2742 4616
rect 2890 4624 2902 4626
rect 2890 4616 2892 4624
rect 2900 4616 2902 4624
rect 2794 4544 2806 4546
rect 2794 4536 2796 4544
rect 2804 4536 2806 4544
rect 2730 3996 2732 4004
rect 2740 3996 2742 4004
rect 2730 3994 2742 3996
rect 2762 4524 2774 4526
rect 2762 4516 2764 4524
rect 2772 4516 2774 4524
rect 2762 3984 2774 4516
rect 2794 4364 2806 4536
rect 2890 4504 2902 4616
rect 3018 4624 3030 4626
rect 3018 4616 3020 4624
rect 3028 4616 3030 4624
rect 2890 4496 2892 4504
rect 2900 4496 2902 4504
rect 2890 4494 2902 4496
rect 2922 4604 2934 4606
rect 2922 4596 2924 4604
rect 2932 4596 2934 4604
rect 2794 4356 2796 4364
rect 2804 4356 2806 4364
rect 2794 4354 2806 4356
rect 2858 4304 2870 4306
rect 2858 4296 2860 4304
rect 2868 4296 2870 4304
rect 2826 4024 2838 4026
rect 2826 4016 2828 4024
rect 2836 4016 2838 4024
rect 2762 3976 2764 3984
rect 2772 3976 2774 3984
rect 2762 3974 2774 3976
rect 2794 3984 2806 3986
rect 2794 3976 2796 3984
rect 2804 3976 2806 3984
rect 2698 3936 2700 3944
rect 2708 3936 2710 3944
rect 2698 3934 2710 3936
rect 2666 3876 2668 3884
rect 2676 3876 2678 3884
rect 2666 3874 2678 3876
rect 2730 3924 2742 3926
rect 2730 3916 2732 3924
rect 2740 3916 2742 3924
rect 2730 3704 2742 3916
rect 2762 3924 2774 3926
rect 2762 3916 2764 3924
rect 2772 3916 2774 3924
rect 2762 3724 2774 3916
rect 2794 3884 2806 3976
rect 2794 3876 2796 3884
rect 2804 3876 2806 3884
rect 2794 3874 2806 3876
rect 2826 3846 2838 4016
rect 2858 4004 2870 4296
rect 2922 4264 2934 4596
rect 3018 4484 3030 4616
rect 3112 4614 3160 4640
rect 3112 4606 3114 4614
rect 3122 4606 3126 4614
rect 3134 4606 3138 4614
rect 3146 4606 3150 4614
rect 3158 4606 3160 4614
rect 3242 4624 3254 4626
rect 3242 4616 3244 4624
rect 3252 4616 3254 4624
rect 3018 4476 3020 4484
rect 3028 4476 3030 4484
rect 3018 4474 3030 4476
rect 3050 4484 3062 4486
rect 3050 4476 3052 4484
rect 3060 4476 3062 4484
rect 2922 4256 2924 4264
rect 2932 4256 2934 4264
rect 2922 4254 2934 4256
rect 2954 4384 2966 4386
rect 2954 4376 2956 4384
rect 2964 4376 2966 4384
rect 2922 4224 2934 4226
rect 2922 4216 2924 4224
rect 2932 4216 2934 4224
rect 2858 3996 2860 4004
rect 2868 3996 2870 4004
rect 2858 3994 2870 3996
rect 2890 4084 2902 4086
rect 2890 4076 2892 4084
rect 2900 4076 2902 4084
rect 2858 3964 2870 3966
rect 2858 3956 2860 3964
rect 2868 3956 2870 3964
rect 2858 3924 2870 3956
rect 2858 3916 2860 3924
rect 2868 3916 2870 3924
rect 2858 3914 2870 3916
rect 2890 3864 2902 4076
rect 2890 3856 2892 3864
rect 2900 3856 2902 3864
rect 2890 3854 2902 3856
rect 2762 3716 2764 3724
rect 2772 3716 2774 3724
rect 2762 3714 2774 3716
rect 2794 3834 2838 3846
rect 2730 3696 2732 3704
rect 2740 3696 2742 3704
rect 2730 3694 2742 3696
rect 2762 3664 2774 3666
rect 2762 3656 2764 3664
rect 2772 3656 2774 3664
rect 2634 3476 2636 3484
rect 2644 3476 2646 3484
rect 2634 3474 2646 3476
rect 2666 3624 2678 3626
rect 2666 3616 2668 3624
rect 2676 3616 2678 3624
rect 2634 3384 2646 3386
rect 2634 3376 2636 3384
rect 2644 3376 2646 3384
rect 2634 3164 2646 3376
rect 2666 3324 2678 3616
rect 2762 3604 2774 3656
rect 2762 3596 2764 3604
rect 2772 3596 2774 3604
rect 2762 3594 2774 3596
rect 2730 3564 2742 3566
rect 2730 3556 2732 3564
rect 2740 3556 2742 3564
rect 2666 3316 2668 3324
rect 2676 3316 2678 3324
rect 2666 3314 2678 3316
rect 2698 3464 2710 3466
rect 2698 3456 2700 3464
rect 2708 3456 2710 3464
rect 2634 3156 2636 3164
rect 2644 3156 2646 3164
rect 2634 3154 2646 3156
rect 2666 3164 2678 3166
rect 2666 3156 2668 3164
rect 2676 3156 2678 3164
rect 2602 3076 2604 3084
rect 2612 3076 2614 3084
rect 2602 3074 2614 3076
rect 2634 3104 2646 3106
rect 2634 3096 2636 3104
rect 2644 3096 2646 3104
rect 2634 3084 2646 3096
rect 2634 3076 2636 3084
rect 2644 3076 2646 3084
rect 2634 3074 2646 3076
rect 2634 3044 2646 3046
rect 2634 3036 2636 3044
rect 2644 3036 2646 3044
rect 2570 2276 2572 2284
rect 2580 2276 2582 2284
rect 2570 2274 2582 2276
rect 2602 3004 2614 3006
rect 2602 2996 2604 3004
rect 2612 2996 2614 3004
rect 2602 2288 2614 2996
rect 2634 2864 2646 3036
rect 2666 2964 2678 3156
rect 2666 2956 2668 2964
rect 2676 2956 2678 2964
rect 2666 2954 2678 2956
rect 2634 2856 2636 2864
rect 2644 2856 2646 2864
rect 2634 2854 2646 2856
rect 2666 2904 2678 2906
rect 2666 2896 2668 2904
rect 2676 2896 2678 2904
rect 2666 2664 2678 2896
rect 2698 2844 2710 3456
rect 2730 3264 2742 3556
rect 2730 3256 2732 3264
rect 2740 3256 2742 3264
rect 2730 3254 2742 3256
rect 2794 3184 2806 3834
rect 2922 3764 2934 4216
rect 2922 3756 2924 3764
rect 2932 3756 2934 3764
rect 2922 3754 2934 3756
rect 2858 3724 2870 3726
rect 2858 3716 2860 3724
rect 2868 3716 2870 3724
rect 2826 3704 2838 3706
rect 2826 3696 2828 3704
rect 2836 3696 2838 3704
rect 2826 3244 2838 3696
rect 2858 3664 2870 3716
rect 2954 3686 2966 4376
rect 3018 4304 3030 4306
rect 3018 4296 3020 4304
rect 3028 4296 3030 4304
rect 2986 4264 2998 4266
rect 2986 4256 2988 4264
rect 2996 4256 2998 4264
rect 2986 4064 2998 4256
rect 3018 4124 3030 4296
rect 3018 4116 3020 4124
rect 3028 4116 3030 4124
rect 3018 4114 3030 4116
rect 2986 4056 2988 4064
rect 2996 4056 2998 4064
rect 2986 4054 2998 4056
rect 2858 3656 2860 3664
rect 2868 3656 2870 3664
rect 2858 3654 2870 3656
rect 2922 3674 2966 3686
rect 2986 3904 2998 3906
rect 2986 3896 2988 3904
rect 2996 3896 2998 3904
rect 2922 3606 2934 3674
rect 2858 3604 2870 3606
rect 2858 3596 2860 3604
rect 2868 3596 2870 3604
rect 2858 3264 2870 3596
rect 2906 3604 2934 3606
rect 2906 3596 2908 3604
rect 2916 3596 2934 3604
rect 2906 3594 2934 3596
rect 2922 3524 2950 3526
rect 2922 3516 2940 3524
rect 2948 3516 2950 3524
rect 2922 3514 2950 3516
rect 2986 3524 2998 3896
rect 3050 3804 3062 4476
rect 3050 3796 3052 3804
rect 3060 3796 3062 3804
rect 3050 3794 3062 3796
rect 3112 4214 3160 4606
rect 3112 4206 3114 4214
rect 3122 4206 3126 4214
rect 3134 4206 3138 4214
rect 3146 4206 3150 4214
rect 3158 4206 3160 4214
rect 3112 3814 3160 4206
rect 3210 4604 3222 4606
rect 3210 4596 3212 4604
rect 3220 4596 3222 4604
rect 3210 3904 3222 4596
rect 3210 3896 3212 3904
rect 3220 3896 3222 3904
rect 3210 3894 3222 3896
rect 3112 3806 3114 3814
rect 3122 3806 3126 3814
rect 3134 3806 3138 3814
rect 3146 3806 3150 3814
rect 3158 3806 3160 3814
rect 2986 3516 2988 3524
rect 2996 3516 2998 3524
rect 2986 3514 2998 3516
rect 3018 3704 3030 3706
rect 3018 3696 3020 3704
rect 3028 3696 3030 3704
rect 2922 3424 2934 3514
rect 2986 3484 2998 3486
rect 2986 3476 2988 3484
rect 2996 3476 2998 3484
rect 2922 3416 2924 3424
rect 2932 3416 2934 3424
rect 2922 3414 2934 3416
rect 2954 3424 2966 3426
rect 2954 3416 2956 3424
rect 2964 3416 2966 3424
rect 2858 3256 2860 3264
rect 2868 3256 2870 3264
rect 2858 3254 2870 3256
rect 2922 3384 2934 3386
rect 2922 3376 2924 3384
rect 2932 3376 2934 3384
rect 2922 3264 2934 3376
rect 2954 3384 2966 3416
rect 2954 3376 2956 3384
rect 2964 3376 2966 3384
rect 2954 3374 2966 3376
rect 2986 3364 2998 3476
rect 2986 3356 2988 3364
rect 2996 3356 2998 3364
rect 2986 3354 2998 3356
rect 2922 3256 2924 3264
rect 2932 3256 2934 3264
rect 2922 3254 2934 3256
rect 2954 3344 2966 3346
rect 2954 3336 2956 3344
rect 2964 3336 2966 3344
rect 2826 3236 2828 3244
rect 2836 3236 2838 3244
rect 2826 3234 2838 3236
rect 2794 3176 2796 3184
rect 2804 3176 2806 3184
rect 2794 3174 2806 3176
rect 2858 3224 2870 3226
rect 2858 3216 2860 3224
rect 2868 3216 2870 3224
rect 2730 3164 2742 3166
rect 2730 3156 2732 3164
rect 2740 3156 2742 3164
rect 2730 3084 2742 3156
rect 2730 3076 2732 3084
rect 2740 3076 2742 3084
rect 2730 3074 2742 3076
rect 2794 3104 2806 3106
rect 2794 3096 2796 3104
rect 2804 3096 2806 3104
rect 2794 3024 2806 3096
rect 2794 3016 2796 3024
rect 2804 3016 2806 3024
rect 2794 3014 2806 3016
rect 2826 3104 2838 3106
rect 2826 3096 2828 3104
rect 2836 3096 2838 3104
rect 2730 3004 2742 3006
rect 2730 2996 2732 3004
rect 2740 2996 2742 3004
rect 2730 2964 2742 2996
rect 2730 2956 2732 2964
rect 2740 2956 2742 2964
rect 2730 2954 2742 2956
rect 2794 2964 2806 2966
rect 2794 2956 2796 2964
rect 2804 2956 2806 2964
rect 2762 2944 2774 2946
rect 2762 2936 2764 2944
rect 2772 2936 2774 2944
rect 2698 2836 2700 2844
rect 2708 2836 2710 2844
rect 2698 2834 2710 2836
rect 2730 2924 2742 2926
rect 2730 2916 2732 2924
rect 2740 2916 2742 2924
rect 2730 2784 2742 2916
rect 2762 2884 2774 2936
rect 2762 2876 2764 2884
rect 2772 2876 2774 2884
rect 2762 2874 2774 2876
rect 2730 2776 2732 2784
rect 2740 2776 2742 2784
rect 2730 2774 2742 2776
rect 2730 2744 2742 2746
rect 2730 2736 2732 2744
rect 2740 2736 2742 2744
rect 2666 2656 2668 2664
rect 2676 2656 2678 2664
rect 2666 2654 2678 2656
rect 2698 2704 2710 2706
rect 2698 2696 2700 2704
rect 2708 2696 2710 2704
rect 2634 2564 2646 2566
rect 2634 2556 2636 2564
rect 2644 2556 2646 2564
rect 2634 2404 2646 2556
rect 2698 2544 2710 2696
rect 2730 2664 2742 2736
rect 2762 2744 2774 2746
rect 2762 2736 2764 2744
rect 2772 2736 2774 2744
rect 2762 2704 2774 2736
rect 2762 2696 2764 2704
rect 2772 2696 2774 2704
rect 2762 2694 2774 2696
rect 2730 2656 2732 2664
rect 2740 2656 2742 2664
rect 2730 2654 2742 2656
rect 2730 2624 2742 2626
rect 2730 2616 2732 2624
rect 2740 2616 2742 2624
rect 2730 2564 2742 2616
rect 2730 2556 2732 2564
rect 2740 2556 2742 2564
rect 2730 2554 2742 2556
rect 2762 2624 2774 2626
rect 2762 2616 2764 2624
rect 2772 2616 2774 2624
rect 2698 2536 2700 2544
rect 2708 2536 2710 2544
rect 2698 2534 2710 2536
rect 2634 2396 2636 2404
rect 2644 2396 2646 2404
rect 2634 2394 2646 2396
rect 2730 2484 2742 2486
rect 2730 2476 2732 2484
rect 2740 2476 2742 2484
rect 2602 2280 2604 2288
rect 2612 2280 2614 2288
rect 2602 2274 2614 2280
rect 2634 2284 2646 2286
rect 2634 2276 2636 2284
rect 2644 2276 2646 2284
rect 2506 2264 2518 2266
rect 2506 2256 2508 2264
rect 2516 2256 2518 2264
rect 2474 2204 2486 2206
rect 2474 2196 2476 2204
rect 2484 2196 2486 2204
rect 2474 2104 2486 2196
rect 2474 2096 2476 2104
rect 2484 2096 2486 2104
rect 2474 2094 2486 2096
rect 2506 2104 2518 2256
rect 2602 2260 2614 2266
rect 2602 2252 2604 2260
rect 2612 2252 2614 2260
rect 2506 2096 2508 2104
rect 2516 2096 2518 2104
rect 2506 2094 2518 2096
rect 2538 2164 2550 2166
rect 2538 2156 2540 2164
rect 2548 2156 2550 2164
rect 2538 2044 2550 2156
rect 2538 2036 2540 2044
rect 2548 2036 2550 2044
rect 2538 2034 2550 2036
rect 2570 2144 2582 2146
rect 2570 2136 2572 2144
rect 2580 2136 2582 2144
rect 2442 1816 2444 1824
rect 2452 1816 2454 1824
rect 2442 1814 2454 1816
rect 2474 2024 2486 2026
rect 2474 2016 2476 2024
rect 2484 2016 2486 2024
rect 2474 1788 2486 2016
rect 2474 1780 2476 1788
rect 2484 1780 2486 1788
rect 2474 1774 2486 1780
rect 2506 2004 2518 2006
rect 2506 1996 2508 2004
rect 2516 1996 2518 2004
rect 2474 1760 2486 1766
rect 2474 1752 2476 1760
rect 2484 1752 2486 1760
rect 2410 1516 2412 1524
rect 2420 1516 2422 1524
rect 2410 1514 2422 1516
rect 2442 1724 2454 1726
rect 2442 1716 2444 1724
rect 2452 1716 2454 1724
rect 2442 1424 2454 1716
rect 2474 1484 2486 1752
rect 2474 1476 2476 1484
rect 2484 1476 2486 1484
rect 2474 1474 2486 1476
rect 2506 1464 2518 1996
rect 2570 1824 2582 2136
rect 2602 2024 2614 2252
rect 2634 2164 2646 2276
rect 2634 2156 2636 2164
rect 2644 2156 2646 2164
rect 2634 2154 2646 2156
rect 2666 2204 2678 2206
rect 2666 2196 2668 2204
rect 2676 2196 2678 2204
rect 2666 2164 2678 2196
rect 2666 2156 2668 2164
rect 2676 2156 2678 2164
rect 2666 2154 2678 2156
rect 2730 2104 2742 2476
rect 2730 2096 2732 2104
rect 2740 2096 2742 2104
rect 2730 2094 2742 2096
rect 2762 2304 2774 2616
rect 2794 2604 2806 2956
rect 2794 2596 2796 2604
rect 2804 2596 2806 2604
rect 2794 2594 2806 2596
rect 2762 2296 2764 2304
rect 2772 2296 2774 2304
rect 2762 2264 2774 2296
rect 2762 2256 2764 2264
rect 2772 2256 2774 2264
rect 2602 2016 2604 2024
rect 2612 2016 2614 2024
rect 2602 2014 2614 2016
rect 2634 2024 2646 2026
rect 2634 2016 2636 2024
rect 2644 2016 2646 2024
rect 2570 1816 2572 1824
rect 2580 1816 2582 1824
rect 2570 1814 2582 1816
rect 2602 1844 2614 1846
rect 2602 1836 2604 1844
rect 2612 1836 2614 1844
rect 2538 1804 2550 1806
rect 2538 1796 2540 1804
rect 2548 1796 2550 1804
rect 2538 1684 2550 1796
rect 2538 1676 2540 1684
rect 2548 1676 2550 1684
rect 2538 1674 2550 1676
rect 2506 1456 2508 1464
rect 2516 1456 2518 1464
rect 2506 1454 2518 1456
rect 2538 1644 2550 1646
rect 2538 1636 2540 1644
rect 2548 1636 2550 1644
rect 2442 1416 2444 1424
rect 2452 1416 2454 1424
rect 2442 1414 2454 1416
rect 2506 1424 2518 1426
rect 2506 1416 2508 1424
rect 2516 1416 2518 1424
rect 2442 1324 2454 1326
rect 2442 1316 2444 1324
rect 2452 1316 2454 1324
rect 2378 1276 2380 1284
rect 2388 1276 2390 1284
rect 2378 1274 2390 1276
rect 2410 1304 2422 1306
rect 2410 1296 2412 1304
rect 2420 1296 2422 1304
rect 2314 1216 2316 1224
rect 2324 1216 2326 1224
rect 2314 1214 2326 1216
rect 2346 1244 2358 1246
rect 2346 1236 2348 1244
rect 2356 1236 2358 1244
rect 2282 1196 2284 1204
rect 2292 1196 2294 1204
rect 2282 1194 2294 1196
rect 2314 1184 2326 1186
rect 2314 1176 2316 1184
rect 2324 1176 2326 1184
rect 2314 1024 2326 1176
rect 2314 1016 2316 1024
rect 2324 1016 2326 1024
rect 2314 1014 2326 1016
rect 2346 1024 2358 1236
rect 2346 1016 2348 1024
rect 2356 1016 2358 1024
rect 2346 1014 2358 1016
rect 2378 1024 2390 1026
rect 2378 1016 2380 1024
rect 2388 1016 2390 1024
rect 2314 984 2326 986
rect 2314 976 2316 984
rect 2324 976 2326 984
rect 2250 896 2252 904
rect 2260 896 2262 904
rect 2250 894 2262 896
rect 2282 964 2294 966
rect 2282 956 2284 964
rect 2292 956 2294 964
rect 2250 864 2262 866
rect 2250 856 2252 864
rect 2260 856 2262 864
rect 2250 764 2262 856
rect 2282 864 2294 956
rect 2314 904 2326 976
rect 2314 896 2316 904
rect 2324 896 2326 904
rect 2314 894 2326 896
rect 2282 856 2284 864
rect 2292 856 2294 864
rect 2282 854 2294 856
rect 2346 844 2358 846
rect 2346 836 2348 844
rect 2356 836 2358 844
rect 2346 824 2358 836
rect 2346 816 2348 824
rect 2356 816 2358 824
rect 2250 756 2252 764
rect 2260 756 2262 764
rect 2250 754 2262 756
rect 2282 804 2310 806
rect 2282 796 2300 804
rect 2308 796 2310 804
rect 2282 794 2310 796
rect 2282 764 2294 794
rect 2282 756 2284 764
rect 2292 756 2294 764
rect 2282 754 2294 756
rect 2218 736 2220 744
rect 2228 736 2230 744
rect 2218 734 2230 736
rect 2314 744 2326 746
rect 2314 736 2316 744
rect 2324 736 2326 744
rect 2122 724 2134 726
rect 2122 716 2124 724
rect 2132 716 2134 724
rect 2122 624 2134 716
rect 2122 616 2124 624
rect 2132 616 2134 624
rect 2122 614 2134 616
rect 2154 724 2166 726
rect 2154 716 2156 724
rect 2164 716 2166 724
rect 2090 556 2092 564
rect 2100 556 2102 564
rect 2090 554 2102 556
rect 2154 504 2166 716
rect 2250 724 2262 726
rect 2250 716 2252 724
rect 2260 716 2262 724
rect 2154 496 2156 504
rect 2164 496 2166 504
rect 2154 494 2166 496
rect 2186 684 2198 686
rect 2186 676 2188 684
rect 2196 676 2198 684
rect 2122 444 2166 446
rect 2122 436 2124 444
rect 2132 436 2166 444
rect 2122 434 2166 436
rect 2154 424 2166 434
rect 2154 416 2156 424
rect 2164 416 2166 424
rect 2154 414 2166 416
rect 2186 366 2198 676
rect 2218 644 2230 646
rect 2218 636 2220 644
rect 2228 636 2230 644
rect 2218 524 2230 636
rect 2250 604 2262 716
rect 2250 596 2252 604
rect 2260 596 2262 604
rect 2250 594 2262 596
rect 2218 516 2220 524
rect 2228 516 2230 524
rect 2218 514 2230 516
rect 2314 464 2326 736
rect 2314 456 2316 464
rect 2324 456 2326 464
rect 2314 454 2326 456
rect 2154 354 2198 366
rect 2154 304 2166 354
rect 2154 296 2156 304
rect 2164 296 2166 304
rect 2154 294 2166 296
rect 2346 304 2358 816
rect 2378 686 2390 1016
rect 2410 1004 2422 1296
rect 2410 996 2412 1004
rect 2420 996 2422 1004
rect 2410 844 2422 996
rect 2442 944 2454 1316
rect 2442 936 2444 944
rect 2452 936 2454 944
rect 2442 934 2454 936
rect 2410 836 2412 844
rect 2420 836 2422 844
rect 2410 834 2422 836
rect 2442 864 2454 866
rect 2442 856 2444 864
rect 2452 856 2454 864
rect 2442 704 2454 856
rect 2506 784 2518 1416
rect 2538 1124 2550 1636
rect 2570 1604 2582 1606
rect 2570 1596 2572 1604
rect 2580 1596 2582 1604
rect 2570 1464 2582 1596
rect 2570 1456 2572 1464
rect 2580 1456 2582 1464
rect 2570 1454 2582 1456
rect 2538 1116 2540 1124
rect 2548 1116 2550 1124
rect 2538 1114 2550 1116
rect 2570 1324 2582 1326
rect 2570 1316 2572 1324
rect 2580 1316 2582 1324
rect 2538 1084 2550 1086
rect 2538 1076 2540 1084
rect 2548 1076 2550 1084
rect 2538 1004 2550 1076
rect 2538 996 2540 1004
rect 2548 996 2550 1004
rect 2538 994 2550 996
rect 2506 776 2508 784
rect 2516 776 2518 784
rect 2506 774 2518 776
rect 2538 904 2550 906
rect 2538 896 2540 904
rect 2548 896 2550 904
rect 2442 696 2444 704
rect 2452 696 2454 704
rect 2442 694 2454 696
rect 2378 684 2422 686
rect 2378 676 2412 684
rect 2420 676 2422 684
rect 2378 674 2422 676
rect 2346 296 2348 304
rect 2356 296 2358 304
rect 2346 294 2358 296
rect 2378 604 2390 606
rect 2378 596 2380 604
rect 2388 596 2390 604
rect 2154 244 2166 246
rect 2154 236 2156 244
rect 2164 236 2166 244
rect 2058 136 2060 144
rect 2068 136 2070 144
rect 2058 134 2070 136
rect 2090 184 2102 186
rect 2090 176 2092 184
rect 2100 176 2102 184
rect 1962 116 1964 124
rect 1972 116 1974 124
rect 1962 114 1974 116
rect 2058 104 2070 106
rect 2058 96 2060 104
rect 2068 96 2070 104
rect 2058 86 2070 96
rect 2090 86 2102 176
rect 2154 144 2166 236
rect 2378 224 2390 596
rect 2410 604 2422 606
rect 2410 596 2412 604
rect 2420 596 2422 604
rect 2410 524 2422 596
rect 2410 516 2412 524
rect 2420 516 2422 524
rect 2410 514 2422 516
rect 2538 484 2550 896
rect 2570 904 2582 1316
rect 2602 1244 2614 1836
rect 2634 1684 2646 2016
rect 2762 2024 2774 2256
rect 2762 2016 2764 2024
rect 2772 2016 2774 2024
rect 2762 2014 2774 2016
rect 2794 2024 2806 2026
rect 2794 2016 2796 2024
rect 2804 2016 2806 2024
rect 2714 1884 2742 1886
rect 2714 1876 2716 1884
rect 2724 1876 2742 1884
rect 2714 1874 2742 1876
rect 2698 1864 2710 1866
rect 2698 1856 2700 1864
rect 2708 1856 2710 1864
rect 2634 1676 2636 1684
rect 2644 1676 2646 1684
rect 2634 1284 2646 1676
rect 2634 1276 2636 1284
rect 2644 1276 2646 1284
rect 2634 1274 2646 1276
rect 2666 1824 2678 1826
rect 2666 1816 2668 1824
rect 2676 1816 2678 1824
rect 2602 1236 2604 1244
rect 2612 1236 2614 1244
rect 2602 1234 2614 1236
rect 2634 1164 2646 1166
rect 2634 1156 2636 1164
rect 2644 1156 2646 1164
rect 2602 1124 2614 1126
rect 2602 1116 2604 1124
rect 2612 1116 2614 1124
rect 2602 1044 2614 1116
rect 2634 1064 2646 1156
rect 2666 1104 2678 1816
rect 2698 1784 2710 1856
rect 2730 1844 2742 1874
rect 2730 1836 2732 1844
rect 2740 1836 2742 1844
rect 2730 1834 2742 1836
rect 2762 1884 2774 1886
rect 2762 1876 2764 1884
rect 2772 1876 2774 1884
rect 2698 1776 2700 1784
rect 2708 1776 2710 1784
rect 2698 1774 2710 1776
rect 2698 1744 2710 1746
rect 2698 1736 2700 1744
rect 2708 1736 2710 1744
rect 2698 1704 2710 1736
rect 2698 1696 2700 1704
rect 2708 1696 2710 1704
rect 2698 1694 2710 1696
rect 2762 1684 2774 1876
rect 2794 1744 2806 2016
rect 2826 1904 2838 3096
rect 2858 2824 2870 3216
rect 2954 3224 2966 3336
rect 2954 3216 2956 3224
rect 2964 3216 2966 3224
rect 2954 3214 2966 3216
rect 2954 3144 2966 3146
rect 2954 3136 2956 3144
rect 2964 3136 2966 3144
rect 2890 3004 2902 3006
rect 2890 2996 2892 3004
rect 2900 2996 2902 3004
rect 2890 2844 2902 2996
rect 2890 2836 2892 2844
rect 2900 2836 2902 2844
rect 2890 2834 2902 2836
rect 2922 3004 2934 3006
rect 2922 2996 2924 3004
rect 2932 2996 2934 3004
rect 2858 2816 2860 2824
rect 2868 2816 2870 2824
rect 2858 2814 2870 2816
rect 2858 2724 2870 2726
rect 2858 2716 2860 2724
rect 2868 2716 2870 2724
rect 2858 2384 2870 2716
rect 2858 2376 2860 2384
rect 2868 2376 2870 2384
rect 2858 2374 2870 2376
rect 2890 2544 2902 2546
rect 2890 2536 2892 2544
rect 2900 2536 2902 2544
rect 2890 2344 2902 2536
rect 2922 2484 2934 2996
rect 2954 3004 2966 3136
rect 2954 2996 2956 3004
rect 2964 2996 2966 3004
rect 2954 2994 2966 2996
rect 2986 3084 2998 3086
rect 2986 3076 2988 3084
rect 2996 3076 2998 3084
rect 2986 3004 2998 3076
rect 3018 3084 3030 3696
rect 3050 3604 3062 3606
rect 3050 3596 3052 3604
rect 3060 3596 3062 3604
rect 3050 3486 3062 3596
rect 3034 3484 3062 3486
rect 3034 3476 3036 3484
rect 3044 3476 3062 3484
rect 3034 3474 3062 3476
rect 3112 3414 3160 3806
rect 3210 3844 3222 3846
rect 3210 3836 3212 3844
rect 3220 3836 3222 3844
rect 3178 3764 3190 3766
rect 3178 3756 3180 3764
rect 3188 3756 3190 3764
rect 3178 3624 3190 3756
rect 3178 3616 3180 3624
rect 3188 3616 3190 3624
rect 3178 3614 3190 3616
rect 3210 3564 3222 3836
rect 3242 3844 3254 4616
rect 3306 4624 3318 4626
rect 3306 4616 3308 4624
rect 3316 4616 3318 4624
rect 3306 4224 3318 4616
rect 3466 4624 3478 4626
rect 3466 4616 3468 4624
rect 3476 4616 3478 4624
rect 3306 4216 3308 4224
rect 3316 4216 3318 4224
rect 3306 4214 3318 4216
rect 3370 4524 3382 4526
rect 3370 4516 3372 4524
rect 3380 4516 3382 4524
rect 3338 4164 3350 4166
rect 3338 4156 3340 4164
rect 3348 4156 3350 4164
rect 3338 4124 3350 4156
rect 3338 4116 3340 4124
rect 3348 4116 3350 4124
rect 3338 4114 3350 4116
rect 3306 4104 3318 4106
rect 3306 4096 3308 4104
rect 3316 4096 3318 4104
rect 3242 3836 3244 3844
rect 3252 3836 3254 3844
rect 3242 3834 3254 3836
rect 3274 4084 3286 4086
rect 3274 4076 3276 4084
rect 3284 4076 3286 4084
rect 3274 3724 3286 4076
rect 3306 3904 3318 4096
rect 3370 3984 3382 4516
rect 3402 4344 3414 4346
rect 3402 4336 3404 4344
rect 3412 4336 3414 4344
rect 3402 4224 3414 4336
rect 3402 4216 3404 4224
rect 3412 4216 3414 4224
rect 3402 4214 3414 4216
rect 3434 4304 3446 4306
rect 3434 4296 3436 4304
rect 3444 4296 3446 4304
rect 3370 3976 3372 3984
rect 3380 3976 3382 3984
rect 3370 3974 3382 3976
rect 3402 4144 3414 4146
rect 3402 4136 3404 4144
rect 3412 4136 3414 4144
rect 3306 3896 3308 3904
rect 3316 3896 3318 3904
rect 3306 3894 3318 3896
rect 3338 3924 3350 3926
rect 3338 3916 3340 3924
rect 3348 3916 3350 3924
rect 3274 3716 3276 3724
rect 3284 3716 3286 3724
rect 3274 3714 3286 3716
rect 3306 3844 3318 3846
rect 3306 3836 3308 3844
rect 3316 3836 3318 3844
rect 3210 3556 3212 3564
rect 3220 3556 3222 3564
rect 3210 3554 3222 3556
rect 3242 3684 3254 3686
rect 3242 3676 3244 3684
rect 3252 3676 3254 3684
rect 3112 3406 3114 3414
rect 3122 3406 3126 3414
rect 3134 3406 3138 3414
rect 3146 3406 3150 3414
rect 3158 3406 3160 3414
rect 3082 3364 3094 3366
rect 3082 3356 3084 3364
rect 3092 3356 3094 3364
rect 3018 3076 3020 3084
rect 3028 3076 3030 3084
rect 3018 3074 3030 3076
rect 3050 3304 3062 3306
rect 3050 3296 3052 3304
rect 3060 3296 3062 3304
rect 2986 2996 2988 3004
rect 2996 2996 2998 3004
rect 2986 2994 2998 2996
rect 3018 3044 3030 3046
rect 3018 3036 3020 3044
rect 3028 3036 3030 3044
rect 2986 2884 2998 2886
rect 2986 2876 2988 2884
rect 2996 2876 2998 2884
rect 2986 2704 2998 2876
rect 3018 2768 3030 3036
rect 3050 2884 3062 3296
rect 3082 3304 3094 3356
rect 3082 3296 3084 3304
rect 3092 3296 3094 3304
rect 3082 3294 3094 3296
rect 3082 3244 3094 3246
rect 3082 3236 3084 3244
rect 3092 3236 3094 3244
rect 3082 3124 3094 3236
rect 3082 3116 3084 3124
rect 3092 3116 3094 3124
rect 3082 3114 3094 3116
rect 3112 3014 3160 3406
rect 3242 3404 3254 3676
rect 3242 3396 3244 3404
rect 3252 3396 3254 3404
rect 3242 3394 3254 3396
rect 3274 3664 3286 3666
rect 3274 3656 3276 3664
rect 3284 3656 3286 3664
rect 3274 3384 3286 3656
rect 3306 3544 3318 3836
rect 3338 3844 3350 3916
rect 3402 3924 3414 4136
rect 3434 3948 3446 4296
rect 3434 3940 3436 3948
rect 3444 3940 3446 3948
rect 3434 3934 3446 3940
rect 3402 3916 3404 3924
rect 3412 3916 3414 3924
rect 3402 3914 3414 3916
rect 3434 3920 3446 3926
rect 3338 3836 3340 3844
rect 3348 3836 3350 3844
rect 3338 3834 3350 3836
rect 3434 3912 3436 3920
rect 3444 3912 3446 3920
rect 3306 3536 3308 3544
rect 3316 3536 3318 3544
rect 3306 3534 3318 3536
rect 3402 3824 3414 3826
rect 3402 3816 3404 3824
rect 3412 3816 3414 3824
rect 3338 3504 3350 3506
rect 3338 3496 3340 3504
rect 3348 3496 3350 3504
rect 3274 3376 3276 3384
rect 3284 3376 3286 3384
rect 3274 3374 3286 3376
rect 3306 3464 3318 3466
rect 3306 3456 3308 3464
rect 3316 3456 3318 3464
rect 3242 3364 3254 3366
rect 3242 3356 3244 3364
rect 3252 3356 3254 3364
rect 3210 3344 3222 3346
rect 3210 3336 3212 3344
rect 3220 3336 3222 3344
rect 3178 3304 3190 3306
rect 3178 3296 3180 3304
rect 3188 3296 3190 3304
rect 3178 3064 3190 3296
rect 3178 3056 3180 3064
rect 3188 3056 3190 3064
rect 3178 3054 3190 3056
rect 3112 3006 3114 3014
rect 3122 3006 3126 3014
rect 3134 3006 3138 3014
rect 3146 3006 3150 3014
rect 3158 3006 3160 3014
rect 3050 2876 3052 2884
rect 3060 2876 3062 2884
rect 3050 2874 3062 2876
rect 3082 2964 3094 2966
rect 3082 2956 3084 2964
rect 3092 2956 3094 2964
rect 3018 2760 3020 2768
rect 3028 2760 3030 2768
rect 3018 2754 3030 2760
rect 3050 2804 3062 2806
rect 3050 2796 3052 2804
rect 3060 2796 3062 2804
rect 2986 2696 2988 2704
rect 2996 2696 2998 2704
rect 2986 2694 2998 2696
rect 3018 2740 3030 2746
rect 3018 2732 3020 2740
rect 3028 2732 3030 2740
rect 2954 2684 2966 2686
rect 2954 2676 2956 2684
rect 2964 2676 2966 2684
rect 2954 2564 2966 2676
rect 2954 2556 2956 2564
rect 2964 2556 2966 2564
rect 2954 2554 2966 2556
rect 2986 2604 2998 2606
rect 2986 2596 2988 2604
rect 2996 2596 2998 2604
rect 2986 2504 2998 2596
rect 2986 2496 2988 2504
rect 2996 2496 2998 2504
rect 2986 2494 2998 2496
rect 2922 2476 2924 2484
rect 2932 2476 2934 2484
rect 2922 2474 2934 2476
rect 2890 2336 2892 2344
rect 2900 2336 2902 2344
rect 2890 2334 2902 2336
rect 2922 2444 2934 2446
rect 2922 2436 2924 2444
rect 2932 2436 2934 2444
rect 2858 2284 2870 2286
rect 2858 2276 2860 2284
rect 2868 2276 2870 2284
rect 2858 2084 2870 2276
rect 2858 2076 2860 2084
rect 2868 2076 2870 2084
rect 2858 2074 2870 2076
rect 2890 2284 2902 2286
rect 2890 2276 2892 2284
rect 2900 2276 2902 2284
rect 2890 2004 2902 2276
rect 2922 2264 2934 2436
rect 3018 2444 3030 2732
rect 3018 2436 3020 2444
rect 3028 2436 3030 2444
rect 3018 2434 3030 2436
rect 3050 2544 3062 2796
rect 3082 2724 3094 2956
rect 3082 2716 3084 2724
rect 3092 2716 3094 2724
rect 3082 2714 3094 2716
rect 3112 2614 3160 3006
rect 3112 2606 3114 2614
rect 3122 2606 3126 2614
rect 3134 2606 3138 2614
rect 3146 2606 3150 2614
rect 3158 2606 3160 2614
rect 3050 2536 3052 2544
rect 3060 2536 3062 2544
rect 2986 2384 2998 2386
rect 2986 2376 2988 2384
rect 2996 2376 2998 2384
rect 2986 2324 2998 2376
rect 3050 2384 3062 2536
rect 3082 2544 3094 2546
rect 3082 2536 3084 2544
rect 3092 2536 3094 2544
rect 3082 2504 3094 2536
rect 3082 2496 3084 2504
rect 3092 2496 3094 2504
rect 3082 2494 3094 2496
rect 3050 2376 3052 2384
rect 3060 2376 3062 2384
rect 3050 2374 3062 2376
rect 2986 2316 2988 2324
rect 2996 2316 2998 2324
rect 2986 2314 2998 2316
rect 3018 2304 3030 2306
rect 3018 2296 3020 2304
rect 3028 2296 3030 2304
rect 2922 2256 2924 2264
rect 2932 2256 2934 2264
rect 2922 2254 2934 2256
rect 2954 2264 2966 2266
rect 2954 2256 2956 2264
rect 2964 2256 2966 2264
rect 2954 2064 2966 2256
rect 2986 2144 2998 2146
rect 2986 2136 2988 2144
rect 2996 2136 2998 2144
rect 2986 2084 2998 2136
rect 2986 2076 2988 2084
rect 2996 2076 2998 2084
rect 2986 2074 2998 2076
rect 2954 2056 2956 2064
rect 2964 2056 2966 2064
rect 2954 2054 2966 2056
rect 3018 2064 3030 2296
rect 3050 2284 3062 2286
rect 3050 2276 3052 2284
rect 3060 2276 3062 2284
rect 3050 2204 3062 2276
rect 3050 2196 3052 2204
rect 3060 2196 3062 2204
rect 3050 2194 3062 2196
rect 3112 2214 3160 2606
rect 3178 2564 3206 2566
rect 3178 2556 3196 2564
rect 3204 2556 3206 2564
rect 3178 2554 3206 2556
rect 3178 2264 3190 2554
rect 3210 2484 3222 3336
rect 3242 3184 3254 3356
rect 3242 3176 3244 3184
rect 3252 3176 3254 3184
rect 3242 3174 3254 3176
rect 3274 3084 3286 3086
rect 3274 3076 3276 3084
rect 3284 3076 3286 3084
rect 3242 3044 3254 3046
rect 3242 3036 3244 3044
rect 3252 3036 3254 3044
rect 3242 2844 3254 3036
rect 3274 2944 3286 3076
rect 3306 3024 3318 3456
rect 3338 3084 3350 3496
rect 3370 3384 3382 3386
rect 3370 3376 3372 3384
rect 3380 3376 3382 3384
rect 3370 3324 3382 3376
rect 3370 3316 3372 3324
rect 3380 3316 3382 3324
rect 3370 3314 3382 3316
rect 3402 3324 3414 3816
rect 3434 3664 3446 3912
rect 3466 3764 3478 4616
rect 4458 4624 4470 4626
rect 4458 4616 4460 4624
rect 4468 4616 4470 4624
rect 3818 4584 3830 4586
rect 3818 4576 3820 4584
rect 3828 4576 3830 4584
rect 3626 4564 3638 4566
rect 3626 4556 3628 4564
rect 3636 4556 3638 4564
rect 3498 4544 3510 4546
rect 3498 4536 3500 4544
rect 3508 4536 3510 4544
rect 3498 4344 3510 4536
rect 3498 4336 3500 4344
rect 3508 4336 3510 4344
rect 3498 4334 3510 4336
rect 3594 4364 3606 4366
rect 3594 4356 3596 4364
rect 3604 4356 3606 4364
rect 3562 4304 3574 4306
rect 3562 4296 3564 4304
rect 3572 4296 3574 4304
rect 3498 4264 3510 4266
rect 3498 4256 3500 4264
rect 3508 4256 3510 4264
rect 3498 3904 3510 4256
rect 3530 4004 3542 4006
rect 3530 3996 3532 4004
rect 3540 3996 3542 4004
rect 3530 3926 3542 3996
rect 3562 3964 3574 4296
rect 3594 4264 3606 4356
rect 3594 4256 3596 4264
rect 3604 4256 3606 4264
rect 3594 4254 3606 4256
rect 3562 3956 3564 3964
rect 3572 3956 3574 3964
rect 3562 3954 3574 3956
rect 3626 4244 3638 4556
rect 3786 4404 3798 4406
rect 3786 4396 3788 4404
rect 3796 4396 3798 4404
rect 3626 4236 3628 4244
rect 3636 4236 3638 4244
rect 3594 3944 3606 3946
rect 3594 3936 3596 3944
rect 3604 3936 3606 3944
rect 3530 3914 3574 3926
rect 3498 3896 3500 3904
rect 3508 3896 3510 3904
rect 3498 3894 3510 3896
rect 3562 3884 3574 3914
rect 3562 3876 3564 3884
rect 3572 3876 3574 3884
rect 3562 3874 3574 3876
rect 3466 3756 3468 3764
rect 3476 3756 3478 3764
rect 3466 3754 3478 3756
rect 3530 3764 3542 3766
rect 3530 3756 3532 3764
rect 3540 3756 3542 3764
rect 3434 3656 3436 3664
rect 3444 3656 3446 3664
rect 3434 3654 3446 3656
rect 3402 3316 3404 3324
rect 3412 3316 3414 3324
rect 3402 3314 3414 3316
rect 3434 3624 3446 3626
rect 3434 3616 3436 3624
rect 3444 3616 3446 3624
rect 3434 3246 3446 3616
rect 3466 3484 3478 3486
rect 3466 3476 3468 3484
rect 3476 3476 3478 3484
rect 3466 3344 3478 3476
rect 3466 3336 3468 3344
rect 3476 3336 3478 3344
rect 3466 3334 3478 3336
rect 3498 3384 3510 3386
rect 3498 3376 3500 3384
rect 3508 3376 3510 3384
rect 3418 3244 3446 3246
rect 3418 3236 3420 3244
rect 3428 3236 3446 3244
rect 3418 3234 3446 3236
rect 3338 3076 3340 3084
rect 3348 3076 3350 3084
rect 3338 3074 3350 3076
rect 3370 3224 3382 3226
rect 3370 3216 3372 3224
rect 3380 3216 3382 3224
rect 3306 3016 3308 3024
rect 3316 3016 3318 3024
rect 3306 3014 3318 3016
rect 3370 3044 3382 3216
rect 3402 3224 3414 3226
rect 3402 3216 3404 3224
rect 3412 3216 3414 3224
rect 3402 3164 3414 3216
rect 3402 3156 3404 3164
rect 3412 3156 3414 3164
rect 3402 3154 3414 3156
rect 3434 3184 3446 3186
rect 3434 3176 3436 3184
rect 3444 3176 3446 3184
rect 3370 3036 3372 3044
rect 3380 3036 3382 3044
rect 3338 3004 3350 3006
rect 3338 2996 3340 3004
rect 3348 2996 3350 3004
rect 3274 2936 3276 2944
rect 3284 2936 3286 2944
rect 3274 2934 3286 2936
rect 3306 2944 3318 2946
rect 3306 2936 3308 2944
rect 3316 2936 3318 2944
rect 3242 2836 3244 2844
rect 3252 2836 3254 2844
rect 3242 2834 3254 2836
rect 3274 2904 3286 2906
rect 3274 2896 3276 2904
rect 3284 2896 3286 2904
rect 3274 2744 3286 2896
rect 3274 2736 3276 2744
rect 3284 2736 3286 2744
rect 3274 2734 3286 2736
rect 3306 2744 3318 2936
rect 3306 2736 3308 2744
rect 3316 2736 3318 2744
rect 3306 2734 3318 2736
rect 3242 2724 3254 2726
rect 3242 2716 3244 2724
rect 3252 2716 3254 2724
rect 3242 2544 3254 2716
rect 3242 2536 3244 2544
rect 3252 2536 3254 2544
rect 3242 2534 3254 2536
rect 3274 2664 3286 2666
rect 3274 2656 3276 2664
rect 3284 2656 3286 2664
rect 3210 2476 3212 2484
rect 3220 2476 3222 2484
rect 3210 2474 3222 2476
rect 3274 2464 3286 2656
rect 3274 2456 3276 2464
rect 3284 2456 3286 2464
rect 3274 2454 3286 2456
rect 3306 2644 3318 2646
rect 3306 2636 3308 2644
rect 3316 2636 3318 2644
rect 3306 2444 3318 2636
rect 3306 2436 3308 2444
rect 3316 2436 3318 2444
rect 3306 2434 3318 2436
rect 3242 2424 3254 2426
rect 3242 2416 3244 2424
rect 3252 2416 3254 2424
rect 3194 2404 3222 2406
rect 3194 2396 3196 2404
rect 3204 2396 3222 2404
rect 3194 2394 3222 2396
rect 3178 2256 3180 2264
rect 3188 2256 3190 2264
rect 3178 2254 3190 2256
rect 3112 2206 3114 2214
rect 3122 2206 3126 2214
rect 3134 2206 3138 2214
rect 3146 2206 3150 2214
rect 3158 2206 3160 2214
rect 3018 2056 3020 2064
rect 3028 2056 3030 2064
rect 3018 2054 3030 2056
rect 2890 1996 2892 2004
rect 2900 1996 2902 2004
rect 2890 1994 2902 1996
rect 2922 1964 2934 1966
rect 2922 1956 2924 1964
rect 2932 1956 2934 1964
rect 2922 1928 2934 1956
rect 2922 1920 2924 1928
rect 2932 1920 2934 1928
rect 3018 1964 3030 1966
rect 3018 1956 3020 1964
rect 3028 1956 3030 1964
rect 2922 1914 2934 1920
rect 2954 1924 2966 1926
rect 2954 1916 2956 1924
rect 2964 1916 2966 1924
rect 2826 1896 2828 1904
rect 2836 1896 2838 1904
rect 2826 1894 2838 1896
rect 2922 1900 2934 1906
rect 2922 1892 2924 1900
rect 2932 1892 2934 1900
rect 2794 1736 2796 1744
rect 2804 1736 2806 1744
rect 2794 1734 2806 1736
rect 2890 1884 2902 1886
rect 2890 1876 2892 1884
rect 2900 1876 2902 1884
rect 2890 1704 2902 1876
rect 2890 1696 2892 1704
rect 2900 1696 2902 1704
rect 2890 1694 2902 1696
rect 2762 1676 2764 1684
rect 2772 1676 2774 1684
rect 2762 1674 2774 1676
rect 2826 1684 2838 1686
rect 2826 1676 2828 1684
rect 2836 1676 2838 1684
rect 2698 1664 2710 1666
rect 2698 1656 2700 1664
rect 2708 1656 2710 1664
rect 2698 1484 2710 1656
rect 2794 1624 2806 1626
rect 2794 1616 2796 1624
rect 2804 1616 2806 1624
rect 2698 1476 2700 1484
rect 2708 1476 2710 1484
rect 2698 1324 2710 1476
rect 2698 1316 2700 1324
rect 2708 1316 2710 1324
rect 2698 1314 2710 1316
rect 2730 1544 2742 1546
rect 2730 1536 2732 1544
rect 2740 1536 2742 1544
rect 2730 1204 2742 1536
rect 2762 1544 2774 1546
rect 2762 1536 2764 1544
rect 2772 1536 2774 1544
rect 2762 1464 2774 1536
rect 2794 1504 2806 1616
rect 2794 1496 2796 1504
rect 2804 1496 2806 1504
rect 2794 1494 2806 1496
rect 2762 1456 2764 1464
rect 2772 1456 2774 1464
rect 2762 1454 2774 1456
rect 2794 1464 2806 1466
rect 2794 1456 2796 1464
rect 2804 1456 2806 1464
rect 2730 1196 2732 1204
rect 2740 1196 2742 1204
rect 2730 1194 2742 1196
rect 2762 1324 2774 1326
rect 2762 1316 2764 1324
rect 2772 1316 2774 1324
rect 2666 1096 2668 1104
rect 2676 1096 2678 1104
rect 2666 1094 2678 1096
rect 2698 1184 2710 1186
rect 2698 1176 2700 1184
rect 2708 1176 2710 1184
rect 2634 1056 2636 1064
rect 2644 1056 2646 1064
rect 2634 1054 2646 1056
rect 2602 1036 2604 1044
rect 2612 1036 2614 1044
rect 2602 1034 2614 1036
rect 2570 896 2572 904
rect 2580 896 2582 904
rect 2570 894 2582 896
rect 2602 924 2630 926
rect 2602 916 2620 924
rect 2628 916 2630 924
rect 2602 914 2630 916
rect 2666 924 2678 926
rect 2666 916 2668 924
rect 2676 916 2678 924
rect 2570 724 2582 726
rect 2570 716 2572 724
rect 2580 716 2582 724
rect 2570 646 2582 716
rect 2602 724 2614 914
rect 2602 716 2604 724
rect 2612 716 2614 724
rect 2602 714 2614 716
rect 2634 844 2646 846
rect 2634 836 2636 844
rect 2644 836 2646 844
rect 2634 724 2646 836
rect 2634 716 2636 724
rect 2644 716 2646 724
rect 2634 714 2646 716
rect 2666 684 2678 916
rect 2666 676 2668 684
rect 2676 676 2678 684
rect 2666 674 2678 676
rect 2570 644 2598 646
rect 2570 636 2588 644
rect 2596 636 2598 644
rect 2570 634 2598 636
rect 2666 624 2678 626
rect 2666 616 2668 624
rect 2676 616 2678 624
rect 2666 544 2678 616
rect 2698 624 2710 1176
rect 2762 984 2774 1316
rect 2794 1284 2806 1456
rect 2826 1404 2838 1676
rect 2922 1684 2934 1892
rect 2954 1808 2966 1916
rect 3018 1844 3030 1956
rect 3018 1836 3020 1844
rect 3028 1836 3030 1844
rect 3018 1834 3030 1836
rect 3050 1884 3062 1886
rect 3050 1876 3052 1884
rect 3060 1876 3062 1884
rect 2954 1800 2956 1808
rect 2964 1800 2966 1808
rect 2954 1794 2966 1800
rect 3018 1804 3030 1806
rect 3018 1796 3020 1804
rect 3028 1796 3030 1804
rect 2954 1780 2966 1786
rect 2954 1772 2956 1780
rect 2964 1772 2966 1780
rect 2954 1744 2966 1772
rect 2954 1736 2956 1744
rect 2964 1736 2966 1744
rect 2954 1734 2966 1736
rect 2986 1744 2998 1746
rect 2986 1736 2988 1744
rect 2996 1736 2998 1744
rect 2922 1676 2924 1684
rect 2932 1676 2934 1684
rect 2826 1396 2828 1404
rect 2836 1396 2838 1404
rect 2826 1394 2838 1396
rect 2890 1624 2902 1626
rect 2890 1616 2892 1624
rect 2900 1616 2902 1624
rect 2794 1276 2796 1284
rect 2804 1276 2806 1284
rect 2794 1274 2806 1276
rect 2826 1324 2854 1326
rect 2826 1316 2844 1324
rect 2852 1316 2854 1324
rect 2826 1314 2854 1316
rect 2826 1284 2838 1314
rect 2826 1276 2828 1284
rect 2836 1276 2838 1284
rect 2762 976 2764 984
rect 2772 976 2774 984
rect 2762 974 2774 976
rect 2794 1184 2806 1186
rect 2794 1176 2796 1184
rect 2804 1176 2806 1184
rect 2698 616 2700 624
rect 2708 616 2710 624
rect 2698 614 2710 616
rect 2730 944 2742 946
rect 2730 936 2732 944
rect 2740 936 2742 944
rect 2666 536 2668 544
rect 2676 536 2678 544
rect 2666 534 2678 536
rect 2730 524 2742 936
rect 2730 516 2732 524
rect 2740 516 2742 524
rect 2730 514 2742 516
rect 2762 944 2774 946
rect 2762 936 2764 944
rect 2772 936 2774 944
rect 2762 804 2774 936
rect 2794 924 2806 1176
rect 2826 944 2838 1276
rect 2890 1284 2902 1616
rect 2922 1484 2934 1676
rect 2922 1476 2924 1484
rect 2932 1476 2934 1484
rect 2922 1474 2934 1476
rect 2986 1324 2998 1736
rect 3018 1524 3030 1796
rect 3018 1516 3020 1524
rect 3028 1516 3030 1524
rect 3018 1514 3030 1516
rect 3018 1444 3030 1446
rect 3018 1436 3020 1444
rect 3028 1436 3030 1444
rect 3018 1384 3030 1436
rect 3018 1376 3020 1384
rect 3028 1376 3030 1384
rect 3018 1374 3030 1376
rect 2986 1316 2988 1324
rect 2996 1316 2998 1324
rect 2986 1314 2998 1316
rect 3018 1344 3030 1346
rect 3018 1336 3020 1344
rect 3028 1336 3030 1344
rect 2890 1276 2892 1284
rect 2900 1276 2902 1284
rect 2890 1274 2902 1276
rect 2922 1084 2934 1086
rect 2922 1076 2924 1084
rect 2932 1076 2934 1084
rect 2890 1064 2902 1066
rect 2890 1056 2892 1064
rect 2900 1056 2902 1064
rect 2826 936 2828 944
rect 2836 936 2838 944
rect 2826 934 2838 936
rect 2858 984 2870 986
rect 2858 976 2860 984
rect 2868 976 2870 984
rect 2794 916 2796 924
rect 2804 916 2806 924
rect 2794 914 2806 916
rect 2858 884 2870 976
rect 2858 876 2860 884
rect 2868 876 2870 884
rect 2858 874 2870 876
rect 2762 796 2764 804
rect 2772 796 2774 804
rect 2762 564 2774 796
rect 2826 764 2838 766
rect 2826 756 2828 764
rect 2836 756 2838 764
rect 2826 724 2838 756
rect 2826 716 2828 724
rect 2836 716 2838 724
rect 2826 714 2838 716
rect 2826 684 2838 686
rect 2826 676 2828 684
rect 2836 676 2838 684
rect 2762 556 2764 564
rect 2772 556 2774 564
rect 2538 476 2540 484
rect 2548 476 2550 484
rect 2538 474 2550 476
rect 2634 504 2646 506
rect 2634 496 2636 504
rect 2644 496 2646 504
rect 2474 444 2486 446
rect 2474 436 2476 444
rect 2484 436 2486 444
rect 2410 404 2422 406
rect 2410 396 2412 404
rect 2420 396 2422 404
rect 2410 364 2422 396
rect 2410 356 2412 364
rect 2420 356 2422 364
rect 2410 354 2422 356
rect 2410 304 2422 306
rect 2410 296 2412 304
rect 2420 296 2422 304
rect 2410 246 2422 296
rect 2474 246 2486 436
rect 2506 344 2518 346
rect 2506 336 2508 344
rect 2516 336 2518 344
rect 2506 304 2518 336
rect 2506 296 2508 304
rect 2516 296 2518 304
rect 2506 294 2518 296
rect 2538 344 2550 346
rect 2538 336 2540 344
rect 2548 336 2550 344
rect 2410 234 2486 246
rect 2378 216 2380 224
rect 2388 216 2390 224
rect 2378 214 2390 216
rect 2154 136 2156 144
rect 2164 136 2166 144
rect 2154 134 2166 136
rect 2314 204 2326 206
rect 2314 196 2316 204
rect 2324 196 2326 204
rect 2314 144 2326 196
rect 2314 136 2316 144
rect 2324 136 2326 144
rect 2314 134 2326 136
rect 2058 74 2102 86
rect 2122 124 2150 126
rect 2122 116 2140 124
rect 2148 116 2150 124
rect 2122 114 2150 116
rect 2218 124 2294 126
rect 2218 116 2220 124
rect 2228 116 2294 124
rect 2218 114 2294 116
rect 2538 124 2550 336
rect 2634 324 2646 496
rect 2762 504 2774 556
rect 2762 496 2764 504
rect 2772 496 2774 504
rect 2762 494 2774 496
rect 2794 584 2806 586
rect 2794 576 2796 584
rect 2804 576 2806 584
rect 2794 484 2806 576
rect 2826 504 2838 676
rect 2826 496 2828 504
rect 2836 496 2838 504
rect 2826 494 2838 496
rect 2858 524 2870 526
rect 2858 516 2860 524
rect 2868 516 2870 524
rect 2794 476 2796 484
rect 2804 476 2806 484
rect 2794 474 2806 476
rect 2634 316 2636 324
rect 2644 316 2646 324
rect 2634 314 2646 316
rect 2762 424 2774 426
rect 2762 416 2764 424
rect 2772 416 2774 424
rect 2762 304 2774 416
rect 2762 296 2764 304
rect 2772 296 2774 304
rect 2762 294 2774 296
rect 2794 364 2806 366
rect 2794 356 2796 364
rect 2804 356 2806 364
rect 2538 116 2540 124
rect 2548 116 2550 124
rect 2538 114 2550 116
rect 2602 284 2614 286
rect 2602 276 2604 284
rect 2612 276 2614 284
rect 2122 24 2134 114
rect 2282 86 2294 114
rect 2282 74 2454 86
rect 2490 84 2566 86
rect 2490 76 2492 84
rect 2500 76 2556 84
rect 2564 76 2566 84
rect 2490 74 2566 76
rect 2442 46 2454 74
rect 2442 34 2582 46
rect 2602 44 2614 276
rect 2602 36 2604 44
rect 2612 36 2614 44
rect 2602 34 2614 36
rect 2634 284 2662 286
rect 2634 276 2652 284
rect 2660 276 2662 284
rect 2634 274 2662 276
rect 2698 284 2710 286
rect 2698 276 2700 284
rect 2708 276 2710 284
rect 2122 16 2124 24
rect 2132 16 2134 24
rect 2122 14 2134 16
rect 1576 6 1578 14
rect 1586 6 1590 14
rect 1598 6 1602 14
rect 1610 6 1614 14
rect 1622 6 1624 14
rect 1576 -40 1624 6
rect 2570 6 2582 34
rect 2634 6 2646 274
rect 2666 224 2678 226
rect 2666 216 2668 224
rect 2676 216 2678 224
rect 2666 124 2678 216
rect 2666 116 2668 124
rect 2676 116 2678 124
rect 2666 114 2678 116
rect 2698 24 2710 276
rect 2794 204 2806 356
rect 2826 344 2838 346
rect 2826 336 2828 344
rect 2836 336 2838 344
rect 2826 244 2838 336
rect 2858 324 2870 516
rect 2890 484 2902 1056
rect 2922 904 2934 1076
rect 2922 896 2924 904
rect 2932 896 2934 904
rect 2922 894 2934 896
rect 2986 944 2998 946
rect 2986 936 2988 944
rect 2996 936 2998 944
rect 2922 864 2934 866
rect 2922 856 2924 864
rect 2932 856 2934 864
rect 2922 624 2934 856
rect 2986 784 2998 936
rect 2986 776 2988 784
rect 2996 776 2998 784
rect 2986 774 2998 776
rect 3018 744 3030 1336
rect 3050 1304 3062 1876
rect 3112 1814 3160 2206
rect 3178 2084 3190 2086
rect 3178 2076 3180 2084
rect 3188 2076 3190 2084
rect 3178 1864 3190 2076
rect 3210 2004 3222 2394
rect 3242 2284 3254 2416
rect 3242 2276 3244 2284
rect 3252 2276 3254 2284
rect 3242 2274 3254 2276
rect 3306 2384 3318 2386
rect 3306 2376 3308 2384
rect 3316 2376 3318 2384
rect 3274 2264 3286 2266
rect 3274 2256 3276 2264
rect 3284 2256 3286 2264
rect 3210 1996 3212 2004
rect 3220 1996 3222 2004
rect 3210 1994 3222 1996
rect 3242 2104 3254 2106
rect 3242 2096 3244 2104
rect 3252 2096 3254 2104
rect 3178 1856 3180 1864
rect 3188 1856 3190 1864
rect 3178 1854 3190 1856
rect 3210 1944 3222 1946
rect 3210 1936 3212 1944
rect 3220 1936 3222 1944
rect 3112 1806 3114 1814
rect 3122 1806 3126 1814
rect 3134 1806 3138 1814
rect 3146 1806 3150 1814
rect 3158 1806 3160 1814
rect 3082 1764 3094 1766
rect 3082 1756 3084 1764
rect 3092 1756 3094 1764
rect 3082 1524 3094 1756
rect 3082 1516 3084 1524
rect 3092 1516 3094 1524
rect 3082 1514 3094 1516
rect 3050 1296 3052 1304
rect 3060 1296 3062 1304
rect 3050 1294 3062 1296
rect 3112 1414 3160 1806
rect 3210 1804 3222 1936
rect 3242 1824 3254 2096
rect 3274 1964 3286 2256
rect 3306 2224 3318 2376
rect 3306 2216 3308 2224
rect 3316 2216 3318 2224
rect 3306 2214 3318 2216
rect 3274 1956 3276 1964
rect 3284 1956 3286 1964
rect 3274 1954 3286 1956
rect 3306 2164 3318 2166
rect 3306 2156 3308 2164
rect 3316 2156 3318 2164
rect 3306 1964 3318 2156
rect 3338 2064 3350 2996
rect 3370 2944 3382 3036
rect 3402 3064 3414 3066
rect 3402 3056 3404 3064
rect 3412 3056 3414 3064
rect 3402 3004 3414 3056
rect 3402 2996 3404 3004
rect 3412 2996 3414 3004
rect 3402 2994 3414 2996
rect 3434 3004 3446 3176
rect 3434 2996 3436 3004
rect 3444 2996 3446 3004
rect 3434 2994 3446 2996
rect 3466 3184 3478 3186
rect 3466 3176 3468 3184
rect 3476 3176 3478 3184
rect 3370 2936 3372 2944
rect 3380 2936 3382 2944
rect 3370 2934 3382 2936
rect 3402 2964 3414 2966
rect 3402 2956 3404 2964
rect 3412 2956 3414 2964
rect 3402 2844 3414 2956
rect 3466 2964 3478 3176
rect 3498 3044 3510 3376
rect 3530 3344 3542 3756
rect 3530 3336 3532 3344
rect 3540 3336 3542 3344
rect 3530 3334 3542 3336
rect 3562 3464 3574 3466
rect 3562 3456 3564 3464
rect 3572 3456 3574 3464
rect 3498 3036 3500 3044
rect 3508 3036 3510 3044
rect 3498 3034 3510 3036
rect 3530 3104 3542 3106
rect 3530 3096 3532 3104
rect 3540 3096 3542 3104
rect 3466 2956 3468 2964
rect 3476 2956 3478 2964
rect 3466 2954 3478 2956
rect 3418 2924 3478 2926
rect 3418 2916 3420 2924
rect 3428 2916 3478 2924
rect 3418 2914 3478 2916
rect 3466 2864 3478 2914
rect 3530 2904 3542 3096
rect 3530 2896 3532 2904
rect 3540 2896 3542 2904
rect 3530 2894 3542 2896
rect 3466 2856 3468 2864
rect 3476 2856 3478 2864
rect 3466 2854 3478 2856
rect 3402 2836 3404 2844
rect 3412 2836 3414 2844
rect 3402 2834 3414 2836
rect 3434 2844 3446 2846
rect 3434 2836 3436 2844
rect 3444 2836 3446 2844
rect 3402 2724 3414 2726
rect 3402 2716 3404 2724
rect 3412 2716 3414 2724
rect 3402 2564 3414 2716
rect 3434 2604 3446 2836
rect 3530 2784 3542 2786
rect 3530 2776 3532 2784
rect 3540 2776 3542 2784
rect 3530 2724 3542 2776
rect 3530 2716 3532 2724
rect 3540 2716 3542 2724
rect 3530 2714 3542 2716
rect 3434 2596 3436 2604
rect 3444 2596 3446 2604
rect 3434 2594 3446 2596
rect 3466 2624 3478 2626
rect 3466 2616 3468 2624
rect 3476 2616 3478 2624
rect 3402 2556 3404 2564
rect 3412 2556 3414 2564
rect 3402 2554 3414 2556
rect 3434 2564 3446 2566
rect 3434 2556 3436 2564
rect 3444 2556 3446 2564
rect 3402 2504 3414 2506
rect 3402 2496 3404 2504
rect 3412 2496 3414 2504
rect 3338 2056 3340 2064
rect 3348 2056 3350 2064
rect 3338 2054 3350 2056
rect 3370 2284 3382 2286
rect 3370 2276 3372 2284
rect 3380 2276 3382 2284
rect 3306 1956 3308 1964
rect 3316 1956 3318 1964
rect 3306 1954 3318 1956
rect 3338 2004 3350 2006
rect 3338 1996 3340 2004
rect 3348 1996 3350 2004
rect 3338 1926 3350 1996
rect 3370 2004 3382 2276
rect 3402 2184 3414 2496
rect 3434 2504 3446 2556
rect 3434 2496 3436 2504
rect 3444 2496 3446 2504
rect 3434 2494 3446 2496
rect 3434 2464 3446 2466
rect 3434 2456 3436 2464
rect 3444 2456 3446 2464
rect 3434 2264 3446 2456
rect 3466 2404 3478 2616
rect 3466 2396 3468 2404
rect 3476 2396 3478 2404
rect 3466 2394 3478 2396
rect 3498 2604 3510 2606
rect 3498 2596 3500 2604
rect 3508 2596 3510 2604
rect 3434 2256 3436 2264
rect 3444 2256 3446 2264
rect 3434 2254 3446 2256
rect 3402 2176 3404 2184
rect 3412 2176 3414 2184
rect 3402 2174 3414 2176
rect 3466 2204 3478 2206
rect 3466 2196 3468 2204
rect 3476 2196 3478 2204
rect 3370 1996 3372 2004
rect 3380 1996 3382 2004
rect 3370 1994 3382 1996
rect 3402 2104 3414 2106
rect 3402 2096 3404 2104
rect 3412 2096 3414 2104
rect 3402 2004 3414 2096
rect 3402 1996 3404 2004
rect 3412 1996 3414 2004
rect 3402 1994 3414 1996
rect 3306 1924 3318 1926
rect 3306 1916 3308 1924
rect 3316 1916 3318 1924
rect 3306 1864 3318 1916
rect 3338 1924 3366 1926
rect 3338 1916 3356 1924
rect 3364 1916 3366 1924
rect 3338 1914 3366 1916
rect 3466 1924 3478 2196
rect 3498 2084 3510 2596
rect 3530 2544 3542 2546
rect 3530 2536 3532 2544
rect 3540 2536 3542 2544
rect 3530 2304 3542 2536
rect 3530 2296 3532 2304
rect 3540 2296 3542 2304
rect 3530 2294 3542 2296
rect 3498 2076 3500 2084
rect 3508 2076 3510 2084
rect 3498 2074 3510 2076
rect 3530 2164 3542 2166
rect 3530 2156 3532 2164
rect 3540 2156 3542 2164
rect 3530 2004 3542 2156
rect 3530 1996 3532 2004
rect 3540 1996 3542 2004
rect 3530 1994 3542 1996
rect 3466 1916 3468 1924
rect 3476 1916 3478 1924
rect 3466 1914 3478 1916
rect 3530 1904 3542 1906
rect 3530 1896 3532 1904
rect 3540 1896 3542 1904
rect 3402 1884 3414 1886
rect 3402 1876 3404 1884
rect 3412 1876 3414 1884
rect 3306 1856 3308 1864
rect 3316 1856 3318 1864
rect 3306 1854 3318 1856
rect 3338 1864 3350 1866
rect 3338 1856 3340 1864
rect 3348 1856 3350 1864
rect 3242 1816 3244 1824
rect 3252 1816 3254 1824
rect 3242 1814 3254 1816
rect 3274 1824 3286 1826
rect 3274 1816 3276 1824
rect 3284 1816 3286 1824
rect 3210 1796 3212 1804
rect 3220 1796 3222 1804
rect 3210 1794 3222 1796
rect 3210 1764 3222 1766
rect 3210 1756 3212 1764
rect 3220 1756 3222 1764
rect 3210 1484 3222 1756
rect 3210 1476 3212 1484
rect 3220 1476 3222 1484
rect 3210 1474 3222 1476
rect 3242 1684 3254 1686
rect 3242 1676 3244 1684
rect 3252 1676 3254 1684
rect 3112 1406 3114 1414
rect 3122 1406 3126 1414
rect 3134 1406 3138 1414
rect 3146 1406 3150 1414
rect 3158 1406 3160 1414
rect 3050 1164 3062 1166
rect 3050 1156 3052 1164
rect 3060 1156 3062 1164
rect 3050 1126 3062 1156
rect 3050 1114 3094 1126
rect 3082 1084 3094 1114
rect 3082 1076 3084 1084
rect 3092 1076 3094 1084
rect 3082 1074 3094 1076
rect 3112 1014 3160 1406
rect 3210 1424 3222 1426
rect 3210 1416 3212 1424
rect 3220 1416 3222 1424
rect 3210 1384 3222 1416
rect 3210 1376 3212 1384
rect 3220 1376 3222 1384
rect 3210 1374 3222 1376
rect 3178 1324 3190 1326
rect 3178 1316 3180 1324
rect 3188 1316 3190 1324
rect 3178 1124 3190 1316
rect 3242 1264 3254 1676
rect 3274 1304 3286 1816
rect 3306 1524 3318 1526
rect 3306 1516 3308 1524
rect 3316 1516 3318 1524
rect 3306 1444 3318 1516
rect 3306 1436 3308 1444
rect 3316 1436 3318 1444
rect 3306 1434 3318 1436
rect 3274 1296 3276 1304
rect 3284 1296 3286 1304
rect 3274 1294 3286 1296
rect 3242 1256 3244 1264
rect 3252 1256 3254 1264
rect 3242 1254 3254 1256
rect 3274 1264 3286 1266
rect 3274 1256 3276 1264
rect 3284 1256 3286 1264
rect 3178 1116 3180 1124
rect 3188 1116 3190 1124
rect 3178 1114 3190 1116
rect 3210 1184 3222 1186
rect 3210 1176 3212 1184
rect 3220 1176 3222 1184
rect 3112 1006 3114 1014
rect 3122 1006 3126 1014
rect 3134 1006 3138 1014
rect 3146 1006 3150 1014
rect 3158 1006 3160 1014
rect 3050 944 3062 946
rect 3050 936 3052 944
rect 3060 936 3062 944
rect 3050 804 3062 936
rect 3050 796 3052 804
rect 3060 796 3062 804
rect 3050 794 3062 796
rect 3082 944 3094 946
rect 3082 936 3084 944
rect 3092 936 3094 944
rect 3018 736 3020 744
rect 3028 736 3030 744
rect 3018 734 3030 736
rect 3082 664 3094 936
rect 3082 656 3084 664
rect 3092 656 3094 664
rect 3082 654 3094 656
rect 2922 616 2924 624
rect 2932 616 2934 624
rect 2922 614 2934 616
rect 2954 644 2966 646
rect 2954 636 2956 644
rect 2964 636 2966 644
rect 2954 544 2966 636
rect 2954 536 2956 544
rect 2964 536 2966 544
rect 2954 534 2966 536
rect 3050 644 3062 646
rect 3050 636 3052 644
rect 3060 636 3062 644
rect 2986 524 2998 526
rect 2986 516 2988 524
rect 2996 516 2998 524
rect 2986 486 2998 516
rect 2890 476 2892 484
rect 2900 476 2902 484
rect 2890 474 2902 476
rect 2954 474 2998 486
rect 3018 504 3030 506
rect 3018 496 3020 504
rect 3028 496 3030 504
rect 2922 424 2934 426
rect 2922 416 2924 424
rect 2932 416 2934 424
rect 2858 316 2860 324
rect 2868 316 2870 324
rect 2858 314 2870 316
rect 2890 404 2902 406
rect 2890 396 2892 404
rect 2900 396 2902 404
rect 2826 236 2828 244
rect 2836 236 2838 244
rect 2826 234 2838 236
rect 2890 244 2902 396
rect 2922 304 2934 416
rect 2954 404 2966 474
rect 2954 396 2956 404
rect 2964 396 2966 404
rect 2954 394 2966 396
rect 2986 404 2998 406
rect 2986 396 2988 404
rect 2996 396 2998 404
rect 2922 296 2924 304
rect 2932 296 2934 304
rect 2922 294 2934 296
rect 2954 344 2966 346
rect 2954 336 2956 344
rect 2964 336 2966 344
rect 2890 236 2892 244
rect 2900 236 2902 244
rect 2890 234 2902 236
rect 2794 196 2796 204
rect 2804 196 2806 204
rect 2794 194 2806 196
rect 2890 204 2918 206
rect 2890 196 2908 204
rect 2916 196 2918 204
rect 2890 194 2918 196
rect 2826 164 2838 166
rect 2826 156 2828 164
rect 2836 156 2838 164
rect 2730 114 2806 126
rect 2730 104 2742 114
rect 2730 96 2732 104
rect 2740 96 2742 104
rect 2730 94 2742 96
rect 2794 84 2806 114
rect 2794 76 2796 84
rect 2804 76 2806 84
rect 2794 74 2806 76
rect 2826 84 2838 156
rect 2826 76 2828 84
rect 2836 76 2838 84
rect 2826 74 2838 76
rect 2698 16 2700 24
rect 2708 16 2710 24
rect 2698 14 2710 16
rect 2826 44 2838 46
rect 2826 36 2828 44
rect 2836 36 2838 44
rect 2570 -6 2646 6
rect 2826 -34 2838 36
rect 2890 -34 2902 194
rect 2954 164 2966 336
rect 2986 304 2998 396
rect 3018 404 3030 496
rect 3050 504 3062 636
rect 3050 496 3052 504
rect 3060 496 3062 504
rect 3050 494 3062 496
rect 3112 614 3160 1006
rect 3112 606 3114 614
rect 3122 606 3126 614
rect 3134 606 3138 614
rect 3146 606 3150 614
rect 3158 606 3160 614
rect 3018 396 3020 404
rect 3028 396 3030 404
rect 3018 394 3030 396
rect 2986 296 2988 304
rect 2996 296 2998 304
rect 2986 264 2998 296
rect 2986 256 2988 264
rect 2996 256 2998 264
rect 2986 254 2998 256
rect 2954 156 2956 164
rect 2964 156 2966 164
rect 2954 154 2966 156
rect 3050 224 3062 226
rect 3050 216 3052 224
rect 3060 216 3062 224
rect 3018 124 3030 126
rect 3018 116 3020 124
rect 3028 116 3030 124
rect 3018 86 3030 116
rect 3050 124 3062 216
rect 3050 116 3052 124
rect 3060 116 3062 124
rect 3050 114 3062 116
rect 3112 214 3160 606
rect 3210 904 3222 1176
rect 3242 1064 3254 1066
rect 3242 1056 3244 1064
rect 3252 1056 3254 1064
rect 3242 984 3254 1056
rect 3242 976 3244 984
rect 3252 976 3254 984
rect 3242 974 3254 976
rect 3210 896 3212 904
rect 3220 896 3222 904
rect 3210 564 3222 896
rect 3274 724 3286 1256
rect 3338 1104 3350 1856
rect 3370 1844 3382 1846
rect 3370 1836 3372 1844
rect 3380 1836 3382 1844
rect 3370 1724 3382 1836
rect 3370 1716 3372 1724
rect 3380 1716 3382 1724
rect 3370 1714 3382 1716
rect 3402 1644 3414 1876
rect 3530 1804 3542 1896
rect 3530 1796 3532 1804
rect 3540 1796 3542 1804
rect 3530 1794 3542 1796
rect 3562 1884 3574 3456
rect 3594 3424 3606 3936
rect 3626 3844 3638 4236
rect 3690 4344 3702 4346
rect 3690 4336 3692 4344
rect 3700 4336 3702 4344
rect 3690 4164 3702 4336
rect 3690 4156 3692 4164
rect 3700 4156 3702 4164
rect 3690 4154 3702 4156
rect 3722 4284 3734 4286
rect 3722 4276 3724 4284
rect 3732 4276 3734 4284
rect 3658 4084 3670 4086
rect 3658 4076 3660 4084
rect 3668 4076 3670 4084
rect 3658 4004 3670 4076
rect 3658 3996 3660 4004
rect 3668 3996 3670 4004
rect 3658 3994 3670 3996
rect 3690 4004 3702 4006
rect 3690 3996 3692 4004
rect 3700 3996 3702 4004
rect 3626 3836 3628 3844
rect 3636 3836 3638 3844
rect 3626 3834 3638 3836
rect 3658 3904 3670 3906
rect 3658 3896 3660 3904
rect 3668 3896 3670 3904
rect 3626 3744 3638 3746
rect 3626 3736 3628 3744
rect 3636 3736 3638 3744
rect 3626 3704 3638 3736
rect 3626 3696 3628 3704
rect 3636 3696 3638 3704
rect 3626 3694 3638 3696
rect 3658 3624 3670 3896
rect 3690 3884 3702 3996
rect 3690 3876 3692 3884
rect 3700 3876 3702 3884
rect 3690 3874 3702 3876
rect 3722 3884 3734 4276
rect 3722 3876 3724 3884
rect 3732 3876 3734 3884
rect 3658 3616 3660 3624
rect 3668 3616 3670 3624
rect 3658 3614 3670 3616
rect 3690 3844 3702 3846
rect 3690 3836 3692 3844
rect 3700 3836 3702 3844
rect 3594 3416 3596 3424
rect 3604 3416 3606 3424
rect 3594 3414 3606 3416
rect 3626 3504 3638 3506
rect 3626 3496 3628 3504
rect 3636 3496 3638 3504
rect 3626 3424 3638 3496
rect 3626 3416 3628 3424
rect 3636 3416 3638 3424
rect 3626 3404 3638 3416
rect 3626 3396 3628 3404
rect 3636 3396 3638 3404
rect 3626 3394 3638 3396
rect 3658 3484 3670 3486
rect 3658 3476 3660 3484
rect 3668 3476 3670 3484
rect 3626 3324 3638 3326
rect 3626 3316 3628 3324
rect 3636 3316 3638 3324
rect 3594 3064 3606 3066
rect 3594 3056 3596 3064
rect 3604 3056 3606 3064
rect 3594 2864 3606 3056
rect 3594 2856 3596 2864
rect 3604 2856 3606 2864
rect 3594 2854 3606 2856
rect 3594 2704 3606 2706
rect 3594 2696 3596 2704
rect 3604 2696 3606 2704
rect 3594 2584 3606 2696
rect 3626 2704 3638 3316
rect 3658 3084 3670 3476
rect 3690 3364 3702 3836
rect 3690 3356 3692 3364
rect 3700 3356 3702 3364
rect 3690 3354 3702 3356
rect 3658 3076 3660 3084
rect 3668 3076 3670 3084
rect 3658 3074 3670 3076
rect 3690 3164 3702 3166
rect 3690 3156 3692 3164
rect 3700 3156 3702 3164
rect 3690 3086 3702 3156
rect 3722 3124 3734 3876
rect 3754 3904 3766 3906
rect 3754 3896 3756 3904
rect 3764 3896 3766 3904
rect 3754 3864 3766 3896
rect 3754 3856 3756 3864
rect 3764 3856 3766 3864
rect 3754 3564 3766 3856
rect 3786 3724 3798 4396
rect 3818 3764 3830 4576
rect 4234 4544 4246 4546
rect 4234 4536 4236 4544
rect 4244 4536 4246 4544
rect 4138 4504 4150 4506
rect 4138 4496 4140 4504
rect 4148 4496 4150 4504
rect 4074 4464 4086 4466
rect 4074 4456 4076 4464
rect 4084 4456 4086 4464
rect 4074 4284 4086 4456
rect 4074 4276 4076 4284
rect 4084 4276 4086 4284
rect 4074 4274 4086 4276
rect 3978 4224 3990 4226
rect 3978 4216 3980 4224
rect 3988 4216 3990 4224
rect 3978 4124 3990 4216
rect 4074 4204 4086 4206
rect 4074 4196 4076 4204
rect 4084 4196 4086 4204
rect 3978 4116 3980 4124
rect 3988 4116 3990 4124
rect 3978 4114 3990 4116
rect 4010 4184 4022 4186
rect 4010 4176 4012 4184
rect 4020 4176 4022 4184
rect 3978 4084 3990 4086
rect 3978 4076 3980 4084
rect 3988 4076 3990 4084
rect 3978 4006 3990 4076
rect 3882 4004 3990 4006
rect 3882 3996 3884 4004
rect 3892 3996 3990 4004
rect 3882 3994 3990 3996
rect 4010 4004 4022 4176
rect 4010 3996 4012 4004
rect 4020 3996 4022 4004
rect 3946 3964 3958 3966
rect 3946 3956 3948 3964
rect 3956 3956 3958 3964
rect 3850 3904 3862 3906
rect 3850 3896 3852 3904
rect 3860 3896 3862 3904
rect 3850 3844 3862 3896
rect 3850 3836 3852 3844
rect 3860 3836 3862 3844
rect 3850 3834 3862 3836
rect 3818 3756 3820 3764
rect 3828 3756 3830 3764
rect 3818 3754 3830 3756
rect 3786 3716 3788 3724
rect 3796 3716 3798 3724
rect 3786 3714 3798 3716
rect 3850 3684 3862 3686
rect 3850 3676 3852 3684
rect 3860 3676 3862 3684
rect 3754 3556 3756 3564
rect 3764 3556 3766 3564
rect 3754 3554 3766 3556
rect 3818 3604 3830 3606
rect 3818 3596 3820 3604
rect 3828 3596 3830 3604
rect 3818 3564 3830 3596
rect 3818 3556 3820 3564
rect 3828 3556 3830 3564
rect 3818 3554 3830 3556
rect 3850 3504 3862 3676
rect 3850 3496 3852 3504
rect 3860 3496 3862 3504
rect 3850 3494 3862 3496
rect 3946 3504 3958 3956
rect 4010 3944 4022 3996
rect 4010 3936 4012 3944
rect 4020 3936 4022 3944
rect 4010 3934 4022 3936
rect 4074 3944 4086 4196
rect 4138 3984 4150 4496
rect 4202 4324 4214 4326
rect 4202 4316 4204 4324
rect 4212 4316 4214 4324
rect 4202 4184 4214 4316
rect 4202 4176 4204 4184
rect 4212 4176 4214 4184
rect 4202 4174 4214 4176
rect 4202 4144 4214 4146
rect 4202 4136 4204 4144
rect 4212 4136 4214 4144
rect 4138 3976 4140 3984
rect 4148 3976 4150 3984
rect 4138 3974 4150 3976
rect 4170 4004 4182 4006
rect 4170 3996 4172 4004
rect 4180 3996 4182 4004
rect 4074 3936 4076 3944
rect 4084 3936 4086 3944
rect 4074 3934 4086 3936
rect 4138 3944 4150 3946
rect 4138 3936 4140 3944
rect 4148 3936 4150 3944
rect 3978 3924 3990 3926
rect 3978 3916 3980 3924
rect 3988 3916 3990 3924
rect 3978 3704 3990 3916
rect 4106 3924 4118 3926
rect 4106 3916 4108 3924
rect 4116 3916 4118 3924
rect 3978 3696 3980 3704
rect 3988 3696 3990 3704
rect 3978 3524 3990 3696
rect 4010 3764 4022 3766
rect 4010 3756 4012 3764
rect 4020 3756 4022 3764
rect 4010 3704 4022 3756
rect 4106 3744 4118 3916
rect 4138 3864 4150 3936
rect 4170 3924 4182 3996
rect 4170 3916 4172 3924
rect 4180 3916 4182 3924
rect 4170 3914 4182 3916
rect 4138 3856 4140 3864
rect 4148 3856 4150 3864
rect 4138 3854 4150 3856
rect 4106 3736 4108 3744
rect 4116 3736 4118 3744
rect 4106 3734 4118 3736
rect 4170 3804 4182 3806
rect 4170 3796 4172 3804
rect 4180 3796 4182 3804
rect 4010 3696 4012 3704
rect 4020 3696 4022 3704
rect 4010 3564 4022 3696
rect 4010 3556 4012 3564
rect 4020 3556 4022 3564
rect 4010 3554 4022 3556
rect 4042 3724 4054 3726
rect 4042 3716 4044 3724
rect 4052 3716 4054 3724
rect 4042 3604 4054 3716
rect 4042 3596 4044 3604
rect 4052 3596 4054 3604
rect 3978 3516 3980 3524
rect 3988 3516 3990 3524
rect 3978 3514 3990 3516
rect 3946 3496 3948 3504
rect 3956 3496 3958 3504
rect 3946 3494 3958 3496
rect 3754 3484 3766 3486
rect 3754 3476 3756 3484
rect 3764 3476 3766 3484
rect 3754 3444 3766 3476
rect 3754 3436 3756 3444
rect 3764 3436 3766 3444
rect 3754 3434 3766 3436
rect 3786 3464 3798 3466
rect 3786 3456 3788 3464
rect 3796 3456 3798 3464
rect 3786 3406 3798 3456
rect 3914 3444 3926 3446
rect 3914 3436 3916 3444
rect 3924 3436 3926 3444
rect 3786 3394 3862 3406
rect 3850 3366 3862 3394
rect 3722 3116 3724 3124
rect 3732 3116 3734 3124
rect 3722 3114 3734 3116
rect 3754 3364 3766 3366
rect 3754 3356 3756 3364
rect 3764 3356 3766 3364
rect 3690 3084 3718 3086
rect 3690 3076 3708 3084
rect 3716 3076 3718 3084
rect 3690 3074 3718 3076
rect 3658 3004 3670 3006
rect 3658 2996 3660 3004
rect 3668 2996 3670 3004
rect 3658 2884 3670 2996
rect 3658 2876 3660 2884
rect 3668 2876 3670 2884
rect 3658 2874 3670 2876
rect 3690 3004 3702 3006
rect 3690 2996 3692 3004
rect 3700 2996 3702 3004
rect 3626 2696 3628 2704
rect 3636 2696 3638 2704
rect 3626 2694 3638 2696
rect 3658 2664 3670 2666
rect 3658 2656 3660 2664
rect 3668 2656 3670 2664
rect 3594 2576 3596 2584
rect 3604 2576 3606 2584
rect 3594 2574 3606 2576
rect 3626 2604 3638 2606
rect 3626 2596 3628 2604
rect 3636 2596 3638 2604
rect 3626 2304 3638 2596
rect 3626 2296 3628 2304
rect 3636 2296 3638 2304
rect 3626 2294 3638 2296
rect 3594 2284 3606 2286
rect 3594 2276 3596 2284
rect 3604 2276 3606 2284
rect 3594 2004 3606 2276
rect 3594 1996 3596 2004
rect 3604 1996 3606 2004
rect 3594 1994 3606 1996
rect 3626 2244 3638 2246
rect 3626 2236 3628 2244
rect 3636 2236 3638 2244
rect 3626 1966 3638 2236
rect 3658 2084 3670 2656
rect 3690 2464 3702 2996
rect 3690 2456 3692 2464
rect 3700 2456 3702 2464
rect 3690 2454 3702 2456
rect 3722 2944 3734 2946
rect 3722 2936 3724 2944
rect 3732 2936 3734 2944
rect 3722 2924 3734 2936
rect 3722 2916 3724 2924
rect 3732 2916 3734 2924
rect 3722 2664 3734 2916
rect 3754 2784 3766 3356
rect 3850 3354 3894 3366
rect 3818 3344 3830 3346
rect 3818 3336 3820 3344
rect 3828 3336 3830 3344
rect 3818 3164 3830 3336
rect 3882 3344 3894 3354
rect 3882 3336 3884 3344
rect 3892 3336 3894 3344
rect 3882 3334 3894 3336
rect 3850 3324 3862 3326
rect 3850 3316 3852 3324
rect 3860 3316 3862 3324
rect 3850 3244 3862 3316
rect 3914 3324 3926 3436
rect 3914 3316 3916 3324
rect 3924 3316 3926 3324
rect 3914 3314 3926 3316
rect 3946 3444 3958 3446
rect 3946 3436 3948 3444
rect 3956 3436 3958 3444
rect 3850 3236 3852 3244
rect 3860 3236 3862 3244
rect 3850 3234 3862 3236
rect 3818 3156 3820 3164
rect 3828 3156 3830 3164
rect 3818 3154 3830 3156
rect 3914 3124 3926 3126
rect 3914 3116 3916 3124
rect 3924 3116 3926 3124
rect 3786 3084 3798 3086
rect 3786 3076 3788 3084
rect 3796 3076 3798 3084
rect 3786 2804 3798 3076
rect 3882 3084 3894 3086
rect 3882 3076 3884 3084
rect 3892 3076 3894 3084
rect 3786 2796 3788 2804
rect 3796 2796 3798 2804
rect 3786 2794 3798 2796
rect 3850 2984 3862 2986
rect 3850 2976 3852 2984
rect 3860 2976 3862 2984
rect 3754 2776 3756 2784
rect 3764 2776 3766 2784
rect 3754 2774 3766 2776
rect 3722 2656 3724 2664
rect 3732 2656 3734 2664
rect 3658 2076 3660 2084
rect 3668 2076 3670 2084
rect 3658 2074 3670 2076
rect 3690 2284 3702 2286
rect 3690 2276 3692 2284
rect 3700 2276 3702 2284
rect 3562 1876 3564 1884
rect 3572 1876 3574 1884
rect 3498 1744 3510 1746
rect 3498 1736 3500 1744
rect 3508 1736 3510 1744
rect 3402 1636 3404 1644
rect 3412 1636 3414 1644
rect 3402 1634 3414 1636
rect 3466 1724 3478 1726
rect 3466 1716 3468 1724
rect 3476 1716 3478 1724
rect 3466 1584 3478 1716
rect 3466 1576 3468 1584
rect 3476 1576 3478 1584
rect 3466 1574 3478 1576
rect 3370 1504 3382 1506
rect 3370 1496 3372 1504
rect 3380 1496 3382 1504
rect 3370 1464 3382 1496
rect 3370 1456 3372 1464
rect 3380 1456 3382 1464
rect 3370 1454 3382 1456
rect 3402 1484 3414 1486
rect 3402 1476 3404 1484
rect 3412 1476 3414 1484
rect 3402 1424 3414 1476
rect 3466 1484 3478 1486
rect 3466 1476 3468 1484
rect 3476 1476 3478 1484
rect 3402 1416 3404 1424
rect 3412 1416 3414 1424
rect 3402 1414 3414 1416
rect 3434 1444 3446 1446
rect 3434 1436 3436 1444
rect 3444 1436 3446 1444
rect 3370 1344 3382 1346
rect 3370 1336 3372 1344
rect 3380 1336 3382 1344
rect 3370 1304 3382 1336
rect 3434 1344 3446 1436
rect 3434 1336 3436 1344
rect 3444 1336 3446 1344
rect 3434 1334 3446 1336
rect 3370 1296 3372 1304
rect 3380 1296 3382 1304
rect 3370 1294 3382 1296
rect 3466 1304 3478 1476
rect 3498 1324 3510 1736
rect 3530 1604 3542 1606
rect 3530 1596 3532 1604
rect 3540 1596 3542 1604
rect 3530 1464 3542 1596
rect 3562 1544 3574 1876
rect 3562 1536 3564 1544
rect 3572 1536 3574 1544
rect 3562 1534 3574 1536
rect 3594 1954 3638 1966
rect 3658 2024 3670 2026
rect 3658 2016 3660 2024
rect 3668 2016 3670 2024
rect 3530 1456 3532 1464
rect 3540 1456 3542 1464
rect 3530 1454 3542 1456
rect 3498 1316 3500 1324
rect 3508 1316 3510 1324
rect 3498 1314 3510 1316
rect 3530 1384 3542 1386
rect 3530 1376 3532 1384
rect 3540 1376 3542 1384
rect 3466 1296 3468 1304
rect 3476 1296 3478 1304
rect 3466 1294 3478 1296
rect 3498 1284 3510 1286
rect 3498 1276 3500 1284
rect 3508 1276 3510 1284
rect 3402 1264 3414 1266
rect 3402 1256 3404 1264
rect 3412 1256 3414 1264
rect 3338 1096 3340 1104
rect 3348 1096 3350 1104
rect 3338 1094 3350 1096
rect 3370 1144 3382 1146
rect 3370 1136 3372 1144
rect 3380 1136 3382 1144
rect 3338 984 3350 986
rect 3338 976 3340 984
rect 3348 976 3350 984
rect 3306 884 3318 886
rect 3306 876 3308 884
rect 3316 876 3318 884
rect 3306 844 3318 876
rect 3306 836 3308 844
rect 3316 836 3318 844
rect 3306 834 3318 836
rect 3338 844 3350 976
rect 3370 964 3382 1136
rect 3370 956 3372 964
rect 3380 956 3382 964
rect 3370 954 3382 956
rect 3338 836 3340 844
rect 3348 836 3350 844
rect 3338 834 3350 836
rect 3338 764 3350 766
rect 3338 756 3340 764
rect 3348 756 3350 764
rect 3274 716 3276 724
rect 3284 716 3286 724
rect 3274 714 3286 716
rect 3306 744 3318 746
rect 3306 736 3308 744
rect 3316 736 3318 744
rect 3306 684 3318 736
rect 3306 676 3308 684
rect 3316 676 3318 684
rect 3306 674 3318 676
rect 3242 664 3254 666
rect 3242 656 3244 664
rect 3252 656 3254 664
rect 3242 624 3254 656
rect 3242 616 3244 624
rect 3252 616 3254 624
rect 3242 614 3254 616
rect 3274 584 3286 586
rect 3274 576 3276 584
rect 3284 576 3286 584
rect 3210 556 3212 564
rect 3220 556 3222 564
rect 3210 554 3222 556
rect 3242 564 3254 566
rect 3242 556 3244 564
rect 3252 556 3254 564
rect 3242 404 3254 556
rect 3274 464 3286 576
rect 3306 564 3318 566
rect 3306 556 3308 564
rect 3316 556 3318 564
rect 3306 486 3318 556
rect 3338 524 3350 756
rect 3338 516 3340 524
rect 3348 516 3350 524
rect 3338 514 3350 516
rect 3370 524 3382 526
rect 3370 516 3372 524
rect 3380 516 3382 524
rect 3370 486 3382 516
rect 3306 474 3382 486
rect 3274 456 3276 464
rect 3284 456 3286 464
rect 3274 454 3286 456
rect 3242 396 3244 404
rect 3252 396 3254 404
rect 3242 394 3254 396
rect 3112 206 3114 214
rect 3122 206 3126 214
rect 3134 206 3138 214
rect 3146 206 3150 214
rect 3158 206 3160 214
rect 3018 74 3094 86
rect 3082 64 3094 74
rect 3082 56 3084 64
rect 3092 56 3094 64
rect 3082 54 3094 56
rect 2826 -46 2902 -34
rect 3112 -40 3160 206
rect 3210 344 3222 346
rect 3210 336 3212 344
rect 3220 336 3222 344
rect 3210 104 3222 336
rect 3322 284 3382 286
rect 3322 276 3324 284
rect 3332 276 3382 284
rect 3322 274 3382 276
rect 3402 284 3414 1256
rect 3498 1004 3510 1276
rect 3530 1124 3542 1376
rect 3594 1264 3606 1954
rect 3658 1944 3670 2016
rect 3658 1936 3660 1944
rect 3668 1936 3670 1944
rect 3658 1934 3670 1936
rect 3626 1844 3638 1846
rect 3626 1836 3628 1844
rect 3636 1836 3638 1844
rect 3626 1364 3638 1836
rect 3690 1844 3702 2276
rect 3690 1836 3692 1844
rect 3700 1836 3702 1844
rect 3690 1834 3702 1836
rect 3690 1804 3702 1806
rect 3690 1796 3692 1804
rect 3700 1796 3702 1804
rect 3658 1564 3670 1566
rect 3658 1556 3660 1564
rect 3668 1556 3670 1564
rect 3658 1424 3670 1556
rect 3658 1416 3660 1424
rect 3668 1416 3670 1424
rect 3658 1414 3670 1416
rect 3626 1356 3628 1364
rect 3636 1356 3638 1364
rect 3626 1354 3638 1356
rect 3658 1364 3670 1366
rect 3658 1356 3660 1364
rect 3668 1356 3670 1364
rect 3658 1284 3670 1356
rect 3658 1276 3660 1284
rect 3668 1276 3670 1284
rect 3658 1274 3670 1276
rect 3594 1256 3596 1264
rect 3604 1256 3606 1264
rect 3594 1254 3606 1256
rect 3530 1116 3532 1124
rect 3540 1116 3542 1124
rect 3530 1114 3542 1116
rect 3562 1104 3574 1106
rect 3562 1096 3564 1104
rect 3572 1096 3574 1104
rect 3498 996 3500 1004
rect 3508 996 3510 1004
rect 3498 924 3510 996
rect 3498 916 3500 924
rect 3508 916 3510 924
rect 3498 914 3510 916
rect 3530 1084 3542 1086
rect 3530 1076 3532 1084
rect 3540 1076 3542 1084
rect 3530 924 3542 1076
rect 3530 916 3532 924
rect 3540 916 3542 924
rect 3530 914 3542 916
rect 3562 924 3574 1096
rect 3690 964 3702 1796
rect 3722 1804 3734 2656
rect 3786 2744 3798 2746
rect 3786 2736 3788 2744
rect 3796 2736 3798 2744
rect 3754 2624 3766 2626
rect 3754 2616 3756 2624
rect 3764 2616 3766 2624
rect 3754 2424 3766 2616
rect 3786 2544 3798 2736
rect 3818 2744 3830 2746
rect 3818 2736 3820 2744
rect 3828 2736 3830 2744
rect 3818 2564 3830 2736
rect 3818 2556 3820 2564
rect 3828 2556 3830 2564
rect 3818 2554 3830 2556
rect 3786 2536 3788 2544
rect 3796 2536 3798 2544
rect 3786 2534 3798 2536
rect 3754 2416 3756 2424
rect 3764 2416 3766 2424
rect 3754 2414 3766 2416
rect 3818 2524 3830 2526
rect 3818 2516 3820 2524
rect 3828 2516 3830 2524
rect 3786 2304 3798 2306
rect 3786 2296 3788 2304
rect 3796 2296 3798 2304
rect 3754 2284 3766 2286
rect 3754 2276 3756 2284
rect 3764 2276 3766 2284
rect 3754 1984 3766 2276
rect 3754 1976 3756 1984
rect 3764 1976 3766 1984
rect 3754 1974 3766 1976
rect 3786 2264 3798 2296
rect 3786 2256 3788 2264
rect 3796 2256 3798 2264
rect 3722 1796 3724 1804
rect 3732 1796 3734 1804
rect 3722 1794 3734 1796
rect 3722 1764 3734 1766
rect 3722 1756 3724 1764
rect 3732 1756 3734 1764
rect 3722 1204 3734 1756
rect 3786 1764 3798 2256
rect 3818 1924 3830 2516
rect 3850 2144 3862 2976
rect 3882 2664 3894 3076
rect 3914 2924 3926 3116
rect 3914 2916 3916 2924
rect 3924 2916 3926 2924
rect 3914 2914 3926 2916
rect 3946 2924 3958 3436
rect 3978 3204 3990 3206
rect 3978 3196 3980 3204
rect 3988 3196 3990 3204
rect 3978 3064 3990 3196
rect 3978 3056 3980 3064
rect 3988 3056 3990 3064
rect 3978 3054 3990 3056
rect 4010 3204 4022 3206
rect 4010 3196 4012 3204
rect 4020 3196 4022 3204
rect 4010 3004 4022 3196
rect 4042 3144 4054 3596
rect 4042 3136 4044 3144
rect 4052 3136 4054 3144
rect 4042 3134 4054 3136
rect 4074 3684 4086 3686
rect 4074 3676 4076 3684
rect 4084 3676 4086 3684
rect 4074 3086 4086 3676
rect 4170 3624 4182 3796
rect 4170 3616 4172 3624
rect 4180 3616 4182 3624
rect 4170 3614 4182 3616
rect 4170 3544 4182 3546
rect 4170 3536 4172 3544
rect 4180 3536 4182 3544
rect 4058 3084 4086 3086
rect 4058 3076 4060 3084
rect 4068 3076 4086 3084
rect 4058 3074 4086 3076
rect 4106 3224 4118 3226
rect 4106 3216 4108 3224
rect 4116 3216 4118 3224
rect 4010 2996 4012 3004
rect 4020 2996 4022 3004
rect 4010 2994 4022 2996
rect 4074 3004 4086 3006
rect 4074 2996 4076 3004
rect 4084 2996 4086 3004
rect 3946 2916 3948 2924
rect 3956 2916 3958 2924
rect 3882 2656 3884 2664
rect 3892 2656 3894 2664
rect 3882 2654 3894 2656
rect 3914 2804 3926 2806
rect 3914 2796 3916 2804
rect 3924 2796 3926 2804
rect 3914 2624 3926 2796
rect 3946 2804 3958 2916
rect 4042 2964 4054 2966
rect 4042 2956 4044 2964
rect 4052 2956 4054 2964
rect 3946 2796 3948 2804
rect 3956 2796 3958 2804
rect 3946 2794 3958 2796
rect 4010 2804 4022 2806
rect 4010 2796 4012 2804
rect 4020 2796 4022 2804
rect 3978 2744 3990 2746
rect 3978 2736 3980 2744
rect 3988 2736 3990 2744
rect 3914 2616 3916 2624
rect 3924 2616 3926 2624
rect 3914 2614 3926 2616
rect 3946 2664 3958 2666
rect 3946 2656 3948 2664
rect 3956 2656 3958 2664
rect 3914 2544 3926 2546
rect 3914 2536 3916 2544
rect 3924 2536 3926 2544
rect 3850 2136 3852 2144
rect 3860 2136 3862 2144
rect 3850 2134 3862 2136
rect 3882 2464 3894 2466
rect 3882 2456 3884 2464
rect 3892 2456 3894 2464
rect 3882 2344 3894 2456
rect 3882 2336 3884 2344
rect 3892 2336 3894 2344
rect 3818 1916 3820 1924
rect 3828 1916 3830 1924
rect 3818 1914 3830 1916
rect 3850 2104 3862 2106
rect 3850 2096 3852 2104
rect 3860 2096 3862 2104
rect 3850 1924 3862 2096
rect 3850 1916 3852 1924
rect 3860 1916 3862 1924
rect 3850 1914 3862 1916
rect 3882 1884 3894 2336
rect 3914 2264 3926 2536
rect 3946 2444 3958 2656
rect 3978 2664 3990 2736
rect 3978 2656 3980 2664
rect 3988 2656 3990 2664
rect 3978 2654 3990 2656
rect 3978 2564 3990 2566
rect 3978 2556 3980 2564
rect 3988 2556 3990 2564
rect 3978 2504 3990 2556
rect 3978 2496 3980 2504
rect 3988 2496 3990 2504
rect 3978 2494 3990 2496
rect 3946 2436 3948 2444
rect 3956 2436 3958 2444
rect 3946 2434 3958 2436
rect 3914 2256 3916 2264
rect 3924 2256 3926 2264
rect 3914 2254 3926 2256
rect 3978 2204 3990 2206
rect 3978 2196 3980 2204
rect 3988 2196 3990 2204
rect 3882 1876 3884 1884
rect 3892 1876 3894 1884
rect 3882 1874 3894 1876
rect 3914 2184 3926 2186
rect 3914 2176 3916 2184
rect 3924 2176 3926 2184
rect 3914 2064 3926 2176
rect 3914 2056 3916 2064
rect 3924 2056 3926 2064
rect 3786 1756 3788 1764
rect 3796 1756 3798 1764
rect 3786 1754 3798 1756
rect 3850 1824 3862 1826
rect 3850 1816 3852 1824
rect 3860 1816 3862 1824
rect 3754 1724 3766 1726
rect 3754 1716 3756 1724
rect 3764 1716 3766 1724
rect 3754 1604 3766 1716
rect 3754 1596 3756 1604
rect 3764 1596 3766 1604
rect 3754 1594 3766 1596
rect 3818 1704 3830 1706
rect 3818 1696 3820 1704
rect 3828 1696 3830 1704
rect 3786 1564 3798 1566
rect 3786 1556 3788 1564
rect 3796 1556 3798 1564
rect 3786 1444 3798 1556
rect 3786 1436 3788 1444
rect 3796 1436 3798 1444
rect 3786 1434 3798 1436
rect 3722 1196 3724 1204
rect 3732 1196 3734 1204
rect 3722 1194 3734 1196
rect 3786 1344 3798 1346
rect 3786 1336 3788 1344
rect 3796 1336 3798 1344
rect 3690 956 3692 964
rect 3700 956 3702 964
rect 3562 916 3564 924
rect 3572 916 3574 924
rect 3562 914 3574 916
rect 3658 944 3670 946
rect 3658 936 3660 944
rect 3668 936 3670 944
rect 3530 864 3542 866
rect 3530 856 3532 864
rect 3540 856 3542 864
rect 3498 844 3510 846
rect 3498 836 3500 844
rect 3508 836 3510 844
rect 3466 744 3478 746
rect 3466 736 3468 744
rect 3476 736 3478 744
rect 3434 704 3446 706
rect 3434 696 3436 704
rect 3444 696 3446 704
rect 3434 624 3446 696
rect 3434 616 3436 624
rect 3444 616 3446 624
rect 3434 614 3446 616
rect 3466 484 3478 736
rect 3498 544 3510 836
rect 3498 536 3500 544
rect 3508 536 3510 544
rect 3498 534 3510 536
rect 3530 544 3542 856
rect 3658 864 3670 936
rect 3658 856 3660 864
rect 3668 856 3670 864
rect 3658 854 3670 856
rect 3626 704 3638 706
rect 3626 696 3628 704
rect 3636 696 3638 704
rect 3626 584 3638 696
rect 3626 576 3628 584
rect 3636 576 3638 584
rect 3626 574 3638 576
rect 3530 536 3532 544
rect 3540 536 3542 544
rect 3530 534 3542 536
rect 3658 564 3670 566
rect 3658 556 3660 564
rect 3668 556 3670 564
rect 3658 526 3670 556
rect 3562 514 3670 526
rect 3466 476 3468 484
rect 3476 476 3478 484
rect 3466 474 3478 476
rect 3498 504 3510 506
rect 3498 496 3500 504
rect 3508 496 3510 504
rect 3402 276 3404 284
rect 3412 276 3414 284
rect 3402 274 3414 276
rect 3434 344 3446 346
rect 3434 336 3436 344
rect 3444 336 3446 344
rect 3434 284 3446 336
rect 3434 276 3436 284
rect 3444 276 3446 284
rect 3434 274 3446 276
rect 3370 246 3382 274
rect 3370 234 3446 246
rect 3242 204 3254 206
rect 3242 196 3244 204
rect 3252 196 3254 204
rect 3242 126 3254 196
rect 3274 184 3286 186
rect 3274 176 3276 184
rect 3284 176 3286 184
rect 3274 166 3286 176
rect 3274 164 3334 166
rect 3274 156 3324 164
rect 3332 156 3334 164
rect 3274 154 3334 156
rect 3242 114 3350 126
rect 3210 96 3212 104
rect 3220 96 3222 104
rect 3210 94 3222 96
rect 3338 104 3350 114
rect 3338 96 3340 104
rect 3348 96 3350 104
rect 3338 94 3350 96
rect 3434 64 3446 234
rect 3498 164 3510 496
rect 3562 344 3574 514
rect 3562 336 3564 344
rect 3572 336 3574 344
rect 3562 334 3574 336
rect 3594 384 3606 386
rect 3594 376 3596 384
rect 3604 376 3606 384
rect 3530 324 3542 326
rect 3530 316 3532 324
rect 3540 316 3542 324
rect 3530 264 3542 316
rect 3530 256 3532 264
rect 3540 256 3542 264
rect 3530 254 3542 256
rect 3562 224 3574 226
rect 3562 216 3564 224
rect 3572 216 3574 224
rect 3498 156 3500 164
rect 3508 156 3510 164
rect 3498 154 3510 156
rect 3530 164 3542 166
rect 3530 156 3532 164
rect 3540 156 3542 164
rect 3530 124 3542 156
rect 3530 116 3532 124
rect 3540 116 3542 124
rect 3530 114 3542 116
rect 3562 124 3574 216
rect 3594 224 3606 376
rect 3690 384 3702 956
rect 3754 1184 3766 1186
rect 3754 1176 3756 1184
rect 3764 1176 3766 1184
rect 3754 664 3766 1176
rect 3754 656 3756 664
rect 3764 656 3766 664
rect 3754 654 3766 656
rect 3754 584 3766 586
rect 3754 576 3756 584
rect 3764 576 3766 584
rect 3722 504 3734 506
rect 3722 496 3724 504
rect 3732 496 3734 504
rect 3722 424 3734 496
rect 3754 444 3766 576
rect 3786 584 3798 1336
rect 3818 1084 3830 1696
rect 3850 1284 3862 1816
rect 3914 1604 3926 2056
rect 3946 2064 3958 2066
rect 3946 2056 3948 2064
rect 3956 2056 3958 2064
rect 3946 1984 3958 2056
rect 3978 2004 3990 2196
rect 3978 1996 3980 2004
rect 3988 1996 3990 2004
rect 3978 1994 3990 1996
rect 3946 1976 3948 1984
rect 3956 1976 3958 1984
rect 3946 1974 3958 1976
rect 3914 1596 3916 1604
rect 3924 1596 3926 1604
rect 3914 1594 3926 1596
rect 3978 1884 3990 1886
rect 3978 1876 3980 1884
rect 3988 1876 3990 1884
rect 3914 1564 3926 1566
rect 3914 1556 3916 1564
rect 3924 1556 3926 1564
rect 3850 1276 3852 1284
rect 3860 1276 3862 1284
rect 3850 1274 3862 1276
rect 3882 1344 3894 1346
rect 3882 1336 3884 1344
rect 3892 1336 3894 1344
rect 3818 1076 3820 1084
rect 3828 1076 3830 1084
rect 3818 1074 3830 1076
rect 3882 904 3894 1336
rect 3914 1304 3926 1556
rect 3978 1384 3990 1876
rect 4010 1766 4022 2796
rect 4042 2584 4054 2956
rect 4074 2804 4086 2996
rect 4074 2796 4076 2804
rect 4084 2796 4086 2804
rect 4074 2794 4086 2796
rect 4106 2704 4118 3216
rect 4138 3164 4150 3166
rect 4138 3156 4140 3164
rect 4148 3156 4150 3164
rect 4138 3024 4150 3156
rect 4170 3124 4182 3536
rect 4170 3116 4172 3124
rect 4180 3116 4182 3124
rect 4170 3114 4182 3116
rect 4202 3044 4214 4136
rect 4234 4144 4246 4536
rect 4234 4136 4236 4144
rect 4244 4136 4246 4144
rect 4234 4134 4246 4136
rect 4266 4304 4278 4306
rect 4266 4296 4268 4304
rect 4276 4296 4278 4304
rect 4234 4064 4246 4066
rect 4234 4056 4236 4064
rect 4244 4056 4246 4064
rect 4234 3724 4246 4056
rect 4266 4064 4278 4296
rect 4298 4304 4310 4306
rect 4298 4296 4300 4304
rect 4308 4296 4310 4304
rect 4298 4144 4310 4296
rect 4394 4204 4406 4206
rect 4394 4196 4396 4204
rect 4404 4196 4406 4204
rect 4298 4136 4300 4144
rect 4308 4136 4310 4144
rect 4298 4134 4310 4136
rect 4362 4164 4374 4166
rect 4362 4156 4364 4164
rect 4372 4156 4374 4164
rect 4266 4056 4268 4064
rect 4276 4056 4278 4064
rect 4266 4054 4278 4056
rect 4298 4084 4310 4086
rect 4298 4076 4300 4084
rect 4308 4076 4310 4084
rect 4234 3716 4236 3724
rect 4244 3716 4246 3724
rect 4234 3714 4246 3716
rect 4266 3784 4278 3786
rect 4266 3776 4268 3784
rect 4276 3776 4278 3784
rect 4234 3624 4246 3626
rect 4234 3616 4236 3624
rect 4244 3616 4246 3624
rect 4234 3224 4246 3616
rect 4266 3484 4278 3776
rect 4266 3476 4268 3484
rect 4276 3476 4278 3484
rect 4266 3474 4278 3476
rect 4234 3216 4236 3224
rect 4244 3216 4246 3224
rect 4234 3214 4246 3216
rect 4266 3304 4278 3306
rect 4266 3296 4268 3304
rect 4276 3296 4278 3304
rect 4202 3036 4204 3044
rect 4212 3036 4214 3044
rect 4202 3034 4214 3036
rect 4138 3016 4140 3024
rect 4148 3016 4150 3024
rect 4138 2864 4150 3016
rect 4138 2856 4140 2864
rect 4148 2856 4150 2864
rect 4138 2854 4150 2856
rect 4234 2944 4246 2946
rect 4234 2936 4236 2944
rect 4244 2936 4246 2944
rect 4106 2696 4108 2704
rect 4116 2696 4118 2704
rect 4106 2694 4118 2696
rect 4170 2684 4182 2686
rect 4170 2676 4172 2684
rect 4180 2676 4182 2684
rect 4170 2624 4182 2676
rect 4170 2616 4172 2624
rect 4180 2616 4182 2624
rect 4170 2614 4182 2616
rect 4042 2576 4044 2584
rect 4052 2576 4054 2584
rect 4042 2574 4054 2576
rect 4106 2564 4118 2566
rect 4106 2556 4108 2564
rect 4116 2556 4118 2564
rect 4074 2524 4086 2526
rect 4074 2516 4076 2524
rect 4084 2516 4086 2524
rect 4042 2504 4054 2506
rect 4042 2496 4044 2504
rect 4052 2496 4054 2504
rect 4042 2404 4054 2496
rect 4042 2396 4044 2404
rect 4052 2396 4054 2404
rect 4042 2044 4054 2396
rect 4042 2036 4044 2044
rect 4052 2036 4054 2044
rect 4042 2034 4054 2036
rect 3994 1764 4022 1766
rect 3994 1756 3996 1764
rect 4004 1756 4022 1764
rect 3994 1754 4022 1756
rect 4042 1904 4054 1906
rect 4042 1896 4044 1904
rect 4052 1896 4054 1904
rect 4042 1624 4054 1896
rect 4042 1616 4044 1624
rect 4052 1616 4054 1624
rect 4042 1614 4054 1616
rect 4010 1584 4022 1586
rect 4010 1576 4012 1584
rect 4020 1576 4022 1584
rect 4010 1566 4022 1576
rect 4010 1554 4054 1566
rect 4042 1484 4054 1554
rect 4042 1476 4044 1484
rect 4052 1476 4054 1484
rect 4042 1474 4054 1476
rect 4074 1404 4086 2516
rect 4106 2244 4118 2556
rect 4138 2524 4150 2526
rect 4138 2516 4140 2524
rect 4148 2516 4150 2524
rect 4138 2444 4150 2516
rect 4138 2436 4140 2444
rect 4148 2436 4150 2444
rect 4138 2434 4150 2436
rect 4170 2524 4182 2526
rect 4170 2516 4172 2524
rect 4180 2516 4182 2524
rect 4106 2236 4108 2244
rect 4116 2236 4118 2244
rect 4106 2104 4118 2236
rect 4106 2096 4108 2104
rect 4116 2096 4118 2104
rect 4106 2094 4118 2096
rect 4138 2284 4150 2286
rect 4138 2276 4140 2284
rect 4148 2276 4150 2284
rect 4138 2004 4150 2276
rect 4170 2184 4182 2516
rect 4170 2176 4172 2184
rect 4180 2176 4182 2184
rect 4170 2174 4182 2176
rect 4202 2304 4214 2306
rect 4202 2296 4204 2304
rect 4212 2296 4214 2304
rect 4138 1996 4140 2004
rect 4148 1996 4150 2004
rect 4138 1994 4150 1996
rect 4170 2044 4182 2046
rect 4170 2036 4172 2044
rect 4180 2036 4182 2044
rect 4138 1924 4150 1926
rect 4138 1916 4140 1924
rect 4148 1916 4150 1924
rect 4138 1864 4150 1916
rect 4138 1856 4140 1864
rect 4148 1856 4150 1864
rect 4138 1854 4150 1856
rect 4074 1396 4076 1404
rect 4084 1396 4086 1404
rect 4074 1394 4086 1396
rect 4106 1704 4118 1706
rect 4106 1696 4108 1704
rect 4116 1696 4118 1704
rect 3978 1376 3980 1384
rect 3988 1376 3990 1384
rect 3978 1374 3990 1376
rect 4106 1384 4118 1696
rect 4170 1704 4182 2036
rect 4202 1904 4214 2296
rect 4234 2264 4246 2936
rect 4266 2704 4278 3296
rect 4298 3084 4310 4076
rect 4362 3964 4374 4156
rect 4394 4104 4406 4196
rect 4394 4096 4396 4104
rect 4404 4096 4406 4104
rect 4394 4094 4406 4096
rect 4362 3956 4364 3964
rect 4372 3956 4374 3964
rect 4362 3954 4374 3956
rect 4426 4004 4438 4006
rect 4426 3996 4428 4004
rect 4436 3996 4438 4004
rect 4394 3684 4406 3686
rect 4394 3676 4396 3684
rect 4404 3676 4406 3684
rect 4298 3076 4300 3084
rect 4308 3076 4310 3084
rect 4298 2904 4310 3076
rect 4298 2896 4300 2904
rect 4308 2896 4310 2904
rect 4298 2894 4310 2896
rect 4330 3184 4342 3186
rect 4330 3176 4332 3184
rect 4340 3176 4342 3184
rect 4266 2696 4268 2704
rect 4276 2696 4278 2704
rect 4266 2694 4278 2696
rect 4298 2804 4310 2806
rect 4298 2796 4300 2804
rect 4308 2796 4310 2804
rect 4266 2504 4278 2506
rect 4266 2496 4268 2504
rect 4276 2496 4278 2504
rect 4266 2384 4278 2496
rect 4266 2376 4268 2384
rect 4276 2376 4278 2384
rect 4266 2374 4278 2376
rect 4234 2256 4236 2264
rect 4244 2256 4246 2264
rect 4234 2254 4246 2256
rect 4298 2204 4310 2796
rect 4330 2504 4342 3176
rect 4362 2964 4374 2966
rect 4362 2956 4364 2964
rect 4372 2956 4374 2964
rect 4362 2924 4374 2956
rect 4362 2916 4364 2924
rect 4372 2916 4374 2924
rect 4362 2914 4374 2916
rect 4394 2604 4406 3676
rect 4426 3024 4438 3996
rect 4458 4004 4470 4616
rect 4664 4414 4712 4640
rect 5194 4604 5206 4606
rect 5194 4596 5196 4604
rect 5204 4596 5206 4604
rect 4664 4406 4666 4414
rect 4674 4406 4678 4414
rect 4686 4406 4690 4414
rect 4698 4406 4702 4414
rect 4710 4406 4712 4414
rect 4458 3996 4460 4004
rect 4468 3996 4470 4004
rect 4458 3994 4470 3996
rect 4490 4304 4502 4306
rect 4490 4296 4492 4304
rect 4500 4296 4502 4304
rect 4458 3924 4470 3926
rect 4458 3916 4460 3924
rect 4468 3916 4470 3924
rect 4458 3524 4470 3916
rect 4458 3516 4460 3524
rect 4468 3516 4470 3524
rect 4458 3514 4470 3516
rect 4490 3324 4502 4296
rect 4586 4224 4598 4226
rect 4586 4216 4588 4224
rect 4596 4216 4598 4224
rect 4554 4064 4566 4066
rect 4554 4056 4556 4064
rect 4564 4056 4566 4064
rect 4554 3724 4566 4056
rect 4586 3984 4598 4216
rect 4586 3976 4588 3984
rect 4596 3976 4598 3984
rect 4586 3974 4598 3976
rect 4618 4024 4630 4026
rect 4618 4016 4620 4024
rect 4628 4016 4630 4024
rect 4554 3716 4556 3724
rect 4564 3716 4566 3724
rect 4554 3714 4566 3716
rect 4586 3724 4598 3726
rect 4586 3716 4588 3724
rect 4596 3716 4598 3724
rect 4586 3464 4598 3716
rect 4618 3684 4630 4016
rect 4618 3676 4620 3684
rect 4628 3676 4630 3684
rect 4618 3674 4630 3676
rect 4664 4014 4712 4406
rect 4664 4006 4666 4014
rect 4674 4006 4678 4014
rect 4686 4006 4690 4014
rect 4698 4006 4702 4014
rect 4710 4006 4712 4014
rect 4586 3456 4588 3464
rect 4596 3456 4598 3464
rect 4586 3454 4598 3456
rect 4664 3614 4712 4006
rect 4906 4444 4918 4446
rect 4906 4436 4908 4444
rect 4916 4436 4918 4444
rect 4664 3606 4666 3614
rect 4674 3606 4678 3614
rect 4686 3606 4690 3614
rect 4698 3606 4702 3614
rect 4710 3606 4712 3614
rect 4490 3316 4492 3324
rect 4500 3316 4502 3324
rect 4490 3314 4502 3316
rect 4664 3214 4712 3606
rect 4778 3984 4790 3986
rect 4778 3976 4780 3984
rect 4788 3976 4790 3984
rect 4778 3504 4790 3976
rect 4906 3764 4918 4436
rect 5162 4444 5174 4446
rect 5162 4436 5164 4444
rect 5172 4436 5174 4444
rect 4906 3756 4908 3764
rect 4916 3756 4918 3764
rect 4906 3754 4918 3756
rect 5034 4164 5046 4166
rect 5034 4156 5036 4164
rect 5044 4156 5046 4164
rect 4778 3496 4780 3504
rect 4788 3496 4790 3504
rect 4778 3494 4790 3496
rect 4664 3206 4666 3214
rect 4674 3206 4678 3214
rect 4686 3206 4690 3214
rect 4698 3206 4702 3214
rect 4710 3206 4712 3214
rect 4426 3016 4428 3024
rect 4436 3016 4438 3024
rect 4426 3014 4438 3016
rect 4522 3044 4534 3046
rect 4522 3036 4524 3044
rect 4532 3036 4534 3044
rect 4522 2764 4534 3036
rect 4522 2756 4524 2764
rect 4532 2756 4534 2764
rect 4522 2754 4534 2756
rect 4586 2924 4598 2926
rect 4586 2916 4588 2924
rect 4596 2916 4598 2924
rect 4490 2744 4502 2746
rect 4490 2736 4492 2744
rect 4500 2736 4502 2744
rect 4490 2684 4502 2736
rect 4490 2676 4492 2684
rect 4500 2676 4502 2684
rect 4490 2674 4502 2676
rect 4394 2596 4396 2604
rect 4404 2596 4406 2604
rect 4394 2594 4406 2596
rect 4490 2604 4502 2606
rect 4490 2596 4492 2604
rect 4500 2596 4502 2604
rect 4330 2496 4332 2504
rect 4340 2496 4342 2504
rect 4330 2494 4342 2496
rect 4426 2504 4438 2506
rect 4426 2496 4428 2504
rect 4436 2496 4438 2504
rect 4362 2464 4374 2466
rect 4362 2456 4364 2464
rect 4372 2456 4374 2464
rect 4298 2196 4300 2204
rect 4308 2196 4310 2204
rect 4298 2194 4310 2196
rect 4330 2344 4342 2346
rect 4330 2336 4332 2344
rect 4340 2336 4342 2344
rect 4234 2184 4246 2186
rect 4234 2176 4236 2184
rect 4244 2176 4246 2184
rect 4234 2044 4246 2176
rect 4234 2036 4236 2044
rect 4244 2036 4246 2044
rect 4234 2034 4246 2036
rect 4266 2164 4278 2166
rect 4266 2156 4268 2164
rect 4276 2156 4278 2164
rect 4202 1896 4204 1904
rect 4212 1896 4214 1904
rect 4202 1894 4214 1896
rect 4170 1696 4172 1704
rect 4180 1696 4182 1704
rect 4170 1694 4182 1696
rect 4202 1804 4214 1806
rect 4202 1796 4204 1804
rect 4212 1796 4214 1804
rect 4202 1564 4214 1796
rect 4266 1744 4278 2156
rect 4330 2144 4342 2336
rect 4362 2204 4374 2456
rect 4362 2196 4364 2204
rect 4372 2196 4374 2204
rect 4362 2194 4374 2196
rect 4330 2136 4332 2144
rect 4340 2136 4342 2144
rect 4330 2134 4342 2136
rect 4394 2144 4406 2146
rect 4394 2136 4396 2144
rect 4404 2136 4406 2144
rect 4266 1736 4268 1744
rect 4276 1736 4278 1744
rect 4266 1724 4278 1736
rect 4266 1716 4268 1724
rect 4276 1716 4278 1724
rect 4266 1714 4278 1716
rect 4298 2104 4310 2106
rect 4298 2096 4300 2104
rect 4308 2096 4310 2104
rect 4298 1704 4310 2096
rect 4362 2044 4374 2046
rect 4362 2036 4364 2044
rect 4372 2036 4374 2044
rect 4330 1804 4342 1806
rect 4330 1796 4332 1804
rect 4340 1796 4342 1804
rect 4330 1744 4342 1796
rect 4330 1736 4332 1744
rect 4340 1736 4342 1744
rect 4330 1734 4342 1736
rect 4298 1696 4300 1704
rect 4308 1696 4310 1704
rect 4298 1694 4310 1696
rect 4266 1624 4278 1626
rect 4266 1616 4268 1624
rect 4276 1616 4278 1624
rect 4202 1556 4204 1564
rect 4212 1556 4214 1564
rect 4202 1554 4214 1556
rect 4234 1604 4246 1606
rect 4234 1596 4236 1604
rect 4244 1596 4246 1604
rect 4202 1444 4214 1446
rect 4202 1436 4204 1444
rect 4212 1436 4214 1444
rect 4106 1376 4108 1384
rect 4116 1376 4118 1384
rect 4106 1374 4118 1376
rect 4138 1424 4150 1426
rect 4138 1416 4140 1424
rect 4148 1416 4150 1424
rect 3914 1296 3916 1304
rect 3924 1296 3926 1304
rect 3914 1294 3926 1296
rect 4074 1364 4086 1366
rect 4074 1356 4076 1364
rect 4084 1356 4086 1364
rect 4074 1144 4086 1356
rect 4106 1344 4118 1346
rect 4106 1336 4108 1344
rect 4116 1336 4118 1344
rect 4106 1164 4118 1336
rect 4138 1344 4150 1416
rect 4138 1336 4140 1344
rect 4148 1336 4150 1344
rect 4138 1334 4150 1336
rect 4106 1156 4108 1164
rect 4116 1156 4118 1164
rect 4106 1154 4118 1156
rect 4074 1136 4076 1144
rect 4084 1136 4086 1144
rect 4074 1134 4086 1136
rect 4170 1104 4182 1106
rect 4170 1096 4172 1104
rect 4180 1096 4182 1104
rect 3882 896 3884 904
rect 3892 896 3894 904
rect 3882 894 3894 896
rect 3914 1044 3926 1046
rect 3914 1036 3916 1044
rect 3924 1036 3926 1044
rect 3786 576 3788 584
rect 3796 576 3798 584
rect 3786 524 3798 576
rect 3786 516 3788 524
rect 3796 516 3798 524
rect 3786 514 3798 516
rect 3818 544 3830 546
rect 3818 536 3820 544
rect 3828 536 3830 544
rect 3754 436 3756 444
rect 3764 436 3766 444
rect 3754 434 3766 436
rect 3722 416 3724 424
rect 3732 416 3734 424
rect 3722 414 3734 416
rect 3690 376 3692 384
rect 3700 376 3702 384
rect 3690 374 3702 376
rect 3722 384 3734 386
rect 3722 376 3724 384
rect 3732 376 3734 384
rect 3658 344 3670 346
rect 3658 336 3660 344
rect 3668 336 3670 344
rect 3626 324 3638 326
rect 3626 316 3628 324
rect 3636 316 3638 324
rect 3626 284 3638 316
rect 3626 276 3628 284
rect 3636 276 3638 284
rect 3626 274 3638 276
rect 3658 264 3670 336
rect 3658 256 3660 264
rect 3668 256 3670 264
rect 3658 254 3670 256
rect 3690 344 3702 346
rect 3690 336 3692 344
rect 3700 336 3702 344
rect 3594 216 3596 224
rect 3604 216 3606 224
rect 3594 214 3606 216
rect 3690 144 3702 336
rect 3722 304 3734 376
rect 3722 296 3724 304
rect 3732 296 3734 304
rect 3722 294 3734 296
rect 3754 364 3766 366
rect 3754 356 3756 364
rect 3764 356 3766 364
rect 3754 246 3766 356
rect 3722 234 3766 246
rect 3722 224 3734 234
rect 3722 216 3724 224
rect 3732 216 3734 224
rect 3722 214 3734 216
rect 3754 204 3766 206
rect 3754 196 3756 204
rect 3764 196 3766 204
rect 3690 136 3692 144
rect 3700 136 3702 144
rect 3690 134 3702 136
rect 3722 144 3734 146
rect 3722 136 3724 144
rect 3732 136 3734 144
rect 3562 116 3564 124
rect 3572 116 3574 124
rect 3562 114 3574 116
rect 3722 86 3734 136
rect 3754 124 3766 196
rect 3818 144 3830 536
rect 3914 524 3926 1036
rect 4010 944 4022 946
rect 4010 936 4012 944
rect 4020 936 4022 944
rect 3978 704 3990 706
rect 3978 696 3980 704
rect 3988 696 3990 704
rect 3914 516 3916 524
rect 3924 516 3926 524
rect 3914 514 3926 516
rect 3946 584 3958 586
rect 3946 576 3948 584
rect 3956 576 3958 584
rect 3850 444 3862 446
rect 3850 436 3852 444
rect 3860 436 3862 444
rect 3850 364 3862 436
rect 3946 444 3958 576
rect 3978 564 3990 696
rect 4010 684 4022 936
rect 4138 924 4150 926
rect 4138 916 4140 924
rect 4148 916 4150 924
rect 4106 904 4118 906
rect 4106 896 4108 904
rect 4116 896 4118 904
rect 4106 844 4118 896
rect 4106 836 4108 844
rect 4116 836 4118 844
rect 4106 834 4118 836
rect 4010 676 4012 684
rect 4020 676 4022 684
rect 4010 674 4022 676
rect 3978 556 3980 564
rect 3988 556 3990 564
rect 3978 554 3990 556
rect 4106 564 4118 566
rect 4106 556 4108 564
rect 4116 556 4118 564
rect 4010 544 4022 546
rect 4010 536 4012 544
rect 4020 536 4022 544
rect 4010 484 4022 536
rect 4010 476 4012 484
rect 4020 476 4022 484
rect 4010 474 4022 476
rect 3946 436 3948 444
rect 3956 436 3958 444
rect 3946 434 3958 436
rect 3850 356 3852 364
rect 3860 356 3862 364
rect 3850 354 3862 356
rect 4010 404 4022 406
rect 4010 396 4012 404
rect 4020 396 4022 404
rect 3850 324 3862 326
rect 3850 316 3852 324
rect 3860 316 3862 324
rect 3850 264 3862 316
rect 3850 256 3852 264
rect 3860 256 3862 264
rect 3850 254 3862 256
rect 3882 284 3942 286
rect 3882 276 3932 284
rect 3940 276 3942 284
rect 3882 274 3942 276
rect 3882 264 3894 274
rect 3882 256 3884 264
rect 3892 256 3894 264
rect 3882 254 3894 256
rect 3818 136 3820 144
rect 3828 136 3830 144
rect 3818 134 3830 136
rect 3754 116 3756 124
rect 3764 116 3766 124
rect 3754 114 3766 116
rect 3882 114 3990 126
rect 3882 104 3894 114
rect 3882 96 3884 104
rect 3892 96 3894 104
rect 3882 94 3894 96
rect 3978 104 3990 114
rect 3978 96 3980 104
rect 3988 96 3990 104
rect 3978 94 3990 96
rect 3434 56 3436 64
rect 3444 56 3446 64
rect 3434 54 3446 56
rect 3658 74 3734 86
rect 3658 64 3670 74
rect 3658 56 3660 64
rect 3668 56 3670 64
rect 3658 54 3670 56
rect 4010 44 4022 396
rect 4042 364 4054 366
rect 4042 356 4044 364
rect 4052 356 4054 364
rect 4042 84 4054 356
rect 4106 284 4118 556
rect 4138 544 4150 916
rect 4138 536 4140 544
rect 4148 536 4150 544
rect 4138 534 4150 536
rect 4170 464 4182 1096
rect 4202 1064 4214 1436
rect 4234 1404 4246 1596
rect 4266 1484 4278 1616
rect 4298 1604 4310 1606
rect 4298 1596 4300 1604
rect 4308 1596 4310 1604
rect 4298 1504 4310 1596
rect 4298 1496 4300 1504
rect 4308 1496 4310 1504
rect 4298 1494 4310 1496
rect 4330 1584 4342 1586
rect 4330 1576 4332 1584
rect 4340 1576 4342 1584
rect 4266 1476 4268 1484
rect 4276 1476 4278 1484
rect 4266 1474 4278 1476
rect 4234 1396 4236 1404
rect 4244 1396 4246 1404
rect 4234 1394 4246 1396
rect 4266 1404 4278 1406
rect 4266 1396 4268 1404
rect 4276 1396 4278 1404
rect 4202 1056 4204 1064
rect 4212 1056 4214 1064
rect 4202 1054 4214 1056
rect 4266 1024 4278 1396
rect 4330 1384 4342 1576
rect 4330 1376 4332 1384
rect 4340 1376 4342 1384
rect 4330 1374 4342 1376
rect 4330 1264 4342 1266
rect 4330 1256 4332 1264
rect 4340 1256 4342 1264
rect 4266 1016 4268 1024
rect 4276 1016 4278 1024
rect 4266 1014 4278 1016
rect 4298 1164 4310 1166
rect 4298 1156 4300 1164
rect 4308 1156 4310 1164
rect 4202 1004 4214 1006
rect 4202 996 4204 1004
rect 4212 996 4214 1004
rect 4202 544 4214 996
rect 4202 536 4204 544
rect 4212 536 4214 544
rect 4202 534 4214 536
rect 4266 964 4278 966
rect 4266 956 4268 964
rect 4276 956 4278 964
rect 4266 544 4278 956
rect 4298 884 4310 1156
rect 4330 1044 4342 1256
rect 4362 1084 4374 2036
rect 4394 1964 4406 2136
rect 4394 1956 4396 1964
rect 4404 1956 4406 1964
rect 4394 1954 4406 1956
rect 4426 1744 4438 2496
rect 4490 2304 4502 2596
rect 4586 2604 4598 2916
rect 4618 2824 4630 2826
rect 4618 2816 4620 2824
rect 4628 2816 4630 2824
rect 4618 2784 4630 2816
rect 4618 2776 4620 2784
rect 4628 2776 4630 2784
rect 4618 2774 4630 2776
rect 4664 2814 4712 3206
rect 4664 2806 4666 2814
rect 4674 2806 4678 2814
rect 4686 2806 4690 2814
rect 4698 2806 4702 2814
rect 4710 2806 4712 2814
rect 4586 2596 4588 2604
rect 4596 2596 4598 2604
rect 4490 2296 4492 2304
rect 4500 2296 4502 2304
rect 4490 2294 4502 2296
rect 4522 2544 4534 2546
rect 4522 2536 4524 2544
rect 4532 2536 4534 2544
rect 4458 2244 4470 2246
rect 4458 2236 4460 2244
rect 4468 2236 4470 2244
rect 4458 2064 4470 2236
rect 4458 2056 4460 2064
rect 4468 2056 4470 2064
rect 4458 2054 4470 2056
rect 4522 1904 4534 2536
rect 4586 2344 4598 2596
rect 4586 2336 4588 2344
rect 4596 2336 4598 2344
rect 4586 2334 4598 2336
rect 4618 2584 4630 2586
rect 4618 2576 4620 2584
rect 4628 2576 4630 2584
rect 4586 2164 4598 2166
rect 4586 2156 4588 2164
rect 4596 2156 4598 2164
rect 4586 2084 4598 2156
rect 4618 2124 4630 2576
rect 4618 2116 4620 2124
rect 4628 2116 4630 2124
rect 4618 2114 4630 2116
rect 4664 2414 4712 2806
rect 4664 2406 4666 2414
rect 4674 2406 4678 2414
rect 4686 2406 4690 2414
rect 4698 2406 4702 2414
rect 4710 2406 4712 2414
rect 4586 2076 4588 2084
rect 4596 2076 4598 2084
rect 4586 2074 4598 2076
rect 4618 2084 4630 2086
rect 4618 2076 4620 2084
rect 4628 2076 4630 2084
rect 4522 1896 4524 1904
rect 4532 1896 4534 1904
rect 4522 1894 4534 1896
rect 4586 1964 4598 1966
rect 4586 1956 4588 1964
rect 4596 1956 4598 1964
rect 4426 1736 4428 1744
rect 4436 1736 4438 1744
rect 4426 1734 4438 1736
rect 4554 1744 4566 1746
rect 4554 1736 4556 1744
rect 4564 1736 4566 1744
rect 4426 1704 4438 1706
rect 4426 1696 4428 1704
rect 4436 1696 4438 1704
rect 4362 1076 4364 1084
rect 4372 1076 4374 1084
rect 4362 1074 4374 1076
rect 4394 1544 4406 1546
rect 4394 1536 4396 1544
rect 4404 1536 4406 1544
rect 4330 1036 4332 1044
rect 4340 1036 4342 1044
rect 4330 1034 4342 1036
rect 4362 1024 4374 1026
rect 4362 1016 4364 1024
rect 4372 1016 4374 1024
rect 4330 1004 4342 1006
rect 4330 996 4332 1004
rect 4340 996 4342 1004
rect 4330 904 4342 996
rect 4330 896 4332 904
rect 4340 896 4342 904
rect 4330 894 4342 896
rect 4298 876 4300 884
rect 4308 876 4310 884
rect 4298 874 4310 876
rect 4330 824 4342 826
rect 4330 816 4332 824
rect 4340 816 4342 824
rect 4298 804 4310 806
rect 4298 796 4300 804
rect 4308 796 4310 804
rect 4298 704 4310 796
rect 4330 724 4342 816
rect 4330 716 4332 724
rect 4340 716 4342 724
rect 4330 714 4342 716
rect 4298 696 4300 704
rect 4308 696 4310 704
rect 4298 694 4310 696
rect 4266 536 4268 544
rect 4276 536 4278 544
rect 4266 534 4278 536
rect 4330 624 4342 626
rect 4330 616 4332 624
rect 4340 616 4342 624
rect 4298 524 4310 526
rect 4298 516 4300 524
rect 4308 516 4310 524
rect 4170 456 4172 464
rect 4180 456 4182 464
rect 4170 454 4182 456
rect 4234 504 4246 506
rect 4234 496 4236 504
rect 4244 496 4246 504
rect 4234 404 4246 496
rect 4234 396 4236 404
rect 4244 396 4246 404
rect 4234 394 4246 396
rect 4266 504 4278 506
rect 4266 496 4268 504
rect 4276 496 4278 504
rect 4234 324 4246 326
rect 4234 316 4236 324
rect 4244 316 4246 324
rect 4202 304 4214 306
rect 4202 296 4204 304
rect 4212 296 4214 304
rect 4106 276 4108 284
rect 4116 276 4118 284
rect 4106 274 4118 276
rect 4138 284 4150 286
rect 4138 276 4140 284
rect 4148 276 4150 284
rect 4074 264 4086 266
rect 4074 256 4076 264
rect 4084 256 4086 264
rect 4074 104 4086 256
rect 4074 96 4076 104
rect 4084 96 4086 104
rect 4074 94 4086 96
rect 4106 184 4118 186
rect 4106 176 4108 184
rect 4116 176 4118 184
rect 4106 104 4118 176
rect 4106 96 4108 104
rect 4116 96 4118 104
rect 4106 94 4118 96
rect 4042 76 4044 84
rect 4052 76 4054 84
rect 4042 74 4054 76
rect 4010 36 4012 44
rect 4020 36 4022 44
rect 4010 34 4022 36
rect 4138 24 4150 276
rect 4202 46 4214 296
rect 4234 244 4246 316
rect 4266 324 4278 496
rect 4266 316 4268 324
rect 4276 316 4278 324
rect 4266 314 4278 316
rect 4234 236 4236 244
rect 4244 236 4246 244
rect 4234 234 4246 236
rect 4298 144 4310 516
rect 4330 164 4342 616
rect 4362 444 4374 1016
rect 4394 804 4406 1536
rect 4426 1164 4438 1696
rect 4490 1704 4502 1706
rect 4490 1696 4492 1704
rect 4500 1696 4502 1704
rect 4490 1584 4502 1696
rect 4490 1576 4492 1584
rect 4500 1576 4502 1584
rect 4490 1574 4502 1576
rect 4554 1564 4566 1736
rect 4586 1604 4598 1956
rect 4618 1904 4630 2076
rect 4618 1896 4620 1904
rect 4628 1896 4630 1904
rect 4618 1894 4630 1896
rect 4664 2014 4712 2406
rect 4938 2584 4950 2586
rect 4938 2576 4940 2584
rect 4948 2576 4950 2584
rect 4874 2184 4886 2186
rect 4874 2176 4876 2184
rect 4884 2176 4886 2184
rect 4842 2124 4854 2126
rect 4842 2116 4844 2124
rect 4852 2116 4854 2124
rect 4664 2006 4666 2014
rect 4674 2006 4678 2014
rect 4686 2006 4690 2014
rect 4698 2006 4702 2014
rect 4710 2006 4712 2014
rect 4586 1596 4588 1604
rect 4596 1596 4598 1604
rect 4586 1594 4598 1596
rect 4618 1844 4630 1846
rect 4618 1836 4620 1844
rect 4628 1836 4630 1844
rect 4554 1556 4556 1564
rect 4564 1556 4566 1564
rect 4554 1554 4566 1556
rect 4586 1564 4598 1566
rect 4586 1556 4588 1564
rect 4596 1556 4598 1564
rect 4458 1544 4470 1546
rect 4458 1536 4460 1544
rect 4468 1536 4470 1544
rect 4458 1508 4470 1536
rect 4458 1500 4460 1508
rect 4468 1500 4470 1508
rect 4458 1494 4470 1500
rect 4458 1480 4470 1486
rect 4458 1472 4460 1480
rect 4468 1472 4470 1480
rect 4458 1224 4470 1472
rect 4522 1484 4534 1486
rect 4522 1476 4524 1484
rect 4532 1476 4534 1484
rect 4458 1216 4460 1224
rect 4468 1216 4470 1224
rect 4458 1214 4470 1216
rect 4490 1384 4502 1386
rect 4490 1376 4492 1384
rect 4500 1376 4502 1384
rect 4490 1224 4502 1376
rect 4522 1304 4534 1476
rect 4586 1464 4598 1556
rect 4586 1456 4588 1464
rect 4596 1456 4598 1464
rect 4586 1454 4598 1456
rect 4522 1296 4524 1304
rect 4532 1296 4534 1304
rect 4522 1294 4534 1296
rect 4554 1444 4566 1446
rect 4554 1436 4556 1444
rect 4564 1436 4566 1444
rect 4554 1284 4566 1436
rect 4618 1404 4630 1836
rect 4618 1396 4620 1404
rect 4628 1396 4630 1404
rect 4618 1394 4630 1396
rect 4664 1614 4712 2006
rect 4778 2044 4790 2046
rect 4778 2036 4780 2044
rect 4788 2036 4790 2044
rect 4778 1844 4790 2036
rect 4842 2044 4854 2116
rect 4842 2036 4844 2044
rect 4852 2036 4854 2044
rect 4842 2034 4854 2036
rect 4842 1924 4854 1926
rect 4842 1916 4844 1924
rect 4852 1916 4854 1924
rect 4842 1864 4854 1916
rect 4874 1904 4886 2176
rect 4938 2124 4950 2576
rect 5034 2204 5046 4156
rect 5162 4104 5174 4436
rect 5162 4096 5164 4104
rect 5172 4096 5174 4104
rect 5162 4094 5174 4096
rect 5162 3344 5174 3346
rect 5162 3336 5164 3344
rect 5172 3336 5174 3344
rect 5162 3304 5174 3336
rect 5162 3296 5164 3304
rect 5172 3296 5174 3304
rect 5162 3084 5174 3296
rect 5194 3184 5206 4596
rect 5834 4584 5846 4586
rect 5834 4576 5836 4584
rect 5844 4576 5846 4584
rect 5594 4564 5718 4566
rect 5594 4556 5596 4564
rect 5604 4556 5718 4564
rect 5594 4554 5718 4556
rect 5482 4544 5494 4546
rect 5482 4536 5484 4544
rect 5492 4536 5494 4544
rect 5418 4524 5430 4526
rect 5418 4516 5420 4524
rect 5428 4516 5430 4524
rect 5354 4384 5366 4386
rect 5354 4376 5356 4384
rect 5364 4376 5366 4384
rect 5258 4164 5270 4166
rect 5258 4156 5260 4164
rect 5268 4156 5270 4164
rect 5226 4024 5238 4026
rect 5226 4016 5228 4024
rect 5236 4016 5238 4024
rect 5226 3924 5238 4016
rect 5226 3916 5228 3924
rect 5236 3916 5238 3924
rect 5226 3914 5238 3916
rect 5258 3904 5270 4156
rect 5258 3896 5260 3904
rect 5268 3896 5270 3904
rect 5226 3884 5238 3886
rect 5226 3876 5228 3884
rect 5236 3876 5238 3884
rect 5226 3624 5238 3876
rect 5226 3616 5228 3624
rect 5236 3616 5238 3624
rect 5226 3614 5238 3616
rect 5194 3176 5196 3184
rect 5204 3176 5206 3184
rect 5194 3174 5206 3176
rect 5226 3544 5238 3546
rect 5226 3536 5228 3544
rect 5236 3536 5238 3544
rect 5162 3076 5164 3084
rect 5172 3076 5174 3084
rect 5162 2904 5174 3076
rect 5162 2896 5164 2904
rect 5172 2896 5174 2904
rect 5162 2894 5174 2896
rect 5194 3064 5206 3066
rect 5194 3056 5196 3064
rect 5204 3056 5206 3064
rect 5194 2664 5206 3056
rect 5226 3004 5238 3536
rect 5226 2996 5228 3004
rect 5236 2996 5238 3004
rect 5226 2994 5238 2996
rect 5258 3284 5270 3896
rect 5290 4124 5302 4126
rect 5290 4116 5292 4124
rect 5300 4116 5302 4124
rect 5290 3824 5302 4116
rect 5354 4024 5366 4376
rect 5386 4384 5398 4386
rect 5386 4376 5388 4384
rect 5396 4376 5398 4384
rect 5386 4244 5398 4376
rect 5418 4284 5430 4516
rect 5418 4276 5420 4284
rect 5428 4276 5430 4284
rect 5418 4274 5430 4276
rect 5482 4324 5494 4536
rect 5578 4544 5590 4546
rect 5578 4536 5580 4544
rect 5588 4536 5590 4544
rect 5482 4316 5484 4324
rect 5492 4316 5494 4324
rect 5482 4284 5494 4316
rect 5482 4276 5484 4284
rect 5492 4276 5494 4284
rect 5386 4236 5388 4244
rect 5396 4236 5398 4244
rect 5386 4234 5398 4236
rect 5354 4016 5356 4024
rect 5364 4016 5366 4024
rect 5354 4014 5366 4016
rect 5418 4204 5430 4206
rect 5418 4196 5420 4204
rect 5428 4196 5430 4204
rect 5386 3944 5398 3946
rect 5386 3936 5388 3944
rect 5396 3936 5398 3944
rect 5290 3816 5292 3824
rect 5300 3816 5302 3824
rect 5290 3814 5302 3816
rect 5354 3864 5366 3866
rect 5354 3856 5356 3864
rect 5364 3856 5366 3864
rect 5322 3744 5334 3746
rect 5322 3736 5324 3744
rect 5332 3736 5334 3744
rect 5258 3276 5260 3284
rect 5268 3276 5270 3284
rect 5226 2964 5238 2966
rect 5226 2956 5228 2964
rect 5236 2956 5238 2964
rect 5226 2864 5238 2956
rect 5258 2924 5270 3276
rect 5258 2916 5260 2924
rect 5268 2916 5270 2924
rect 5258 2914 5270 2916
rect 5290 3704 5302 3706
rect 5290 3696 5292 3704
rect 5300 3696 5302 3704
rect 5290 2944 5302 3696
rect 5322 3704 5334 3736
rect 5322 3696 5324 3704
rect 5332 3696 5334 3704
rect 5322 3694 5334 3696
rect 5322 3644 5334 3646
rect 5322 3636 5324 3644
rect 5332 3636 5334 3644
rect 5322 3304 5334 3636
rect 5354 3384 5366 3856
rect 5354 3376 5356 3384
rect 5364 3376 5366 3384
rect 5354 3374 5366 3376
rect 5322 3296 5324 3304
rect 5332 3296 5334 3304
rect 5322 3294 5334 3296
rect 5354 3264 5366 3266
rect 5354 3256 5356 3264
rect 5364 3256 5366 3264
rect 5290 2936 5292 2944
rect 5300 2936 5302 2944
rect 5226 2856 5228 2864
rect 5236 2856 5238 2864
rect 5226 2854 5238 2856
rect 5194 2656 5196 2664
rect 5204 2656 5206 2664
rect 5194 2654 5206 2656
rect 5258 2544 5270 2546
rect 5258 2536 5260 2544
rect 5268 2536 5270 2544
rect 5258 2424 5270 2536
rect 5290 2504 5302 2936
rect 5322 3064 5334 3066
rect 5322 3056 5324 3064
rect 5332 3056 5334 3064
rect 5322 2864 5334 3056
rect 5322 2856 5324 2864
rect 5332 2856 5334 2864
rect 5322 2854 5334 2856
rect 5290 2496 5292 2504
rect 5300 2496 5302 2504
rect 5290 2494 5302 2496
rect 5322 2784 5334 2786
rect 5322 2776 5324 2784
rect 5332 2776 5334 2784
rect 5322 2624 5334 2776
rect 5322 2616 5324 2624
rect 5332 2616 5334 2624
rect 5258 2416 5260 2424
rect 5268 2416 5270 2424
rect 5258 2414 5270 2416
rect 5322 2344 5334 2616
rect 5354 2544 5366 3256
rect 5386 3264 5398 3936
rect 5418 3524 5430 4196
rect 5418 3516 5420 3524
rect 5428 3516 5430 3524
rect 5418 3514 5430 3516
rect 5450 3804 5462 3806
rect 5450 3796 5452 3804
rect 5460 3796 5462 3804
rect 5386 3256 5388 3264
rect 5396 3256 5398 3264
rect 5386 3254 5398 3256
rect 5418 3464 5430 3466
rect 5418 3456 5420 3464
rect 5428 3456 5430 3464
rect 5386 3204 5398 3206
rect 5386 3196 5388 3204
rect 5396 3196 5398 3204
rect 5386 3024 5398 3196
rect 5418 3064 5430 3456
rect 5450 3364 5462 3796
rect 5482 3764 5494 4276
rect 5482 3756 5484 3764
rect 5492 3756 5494 3764
rect 5482 3754 5494 3756
rect 5514 4344 5526 4346
rect 5514 4336 5516 4344
rect 5524 4336 5526 4344
rect 5450 3356 5452 3364
rect 5460 3356 5462 3364
rect 5450 3354 5462 3356
rect 5482 3524 5494 3526
rect 5482 3516 5484 3524
rect 5492 3516 5494 3524
rect 5418 3056 5420 3064
rect 5428 3056 5430 3064
rect 5418 3054 5430 3056
rect 5482 3064 5494 3516
rect 5514 3324 5526 4336
rect 5578 4324 5590 4536
rect 5706 4524 5718 4554
rect 5770 4544 5782 4546
rect 5770 4536 5772 4544
rect 5780 4536 5782 4544
rect 5770 4526 5782 4536
rect 5706 4516 5708 4524
rect 5716 4516 5718 4524
rect 5706 4514 5718 4516
rect 5738 4524 5782 4526
rect 5738 4516 5740 4524
rect 5748 4516 5782 4524
rect 5738 4514 5782 4516
rect 5578 4316 5580 4324
rect 5588 4316 5590 4324
rect 5578 4314 5590 4316
rect 5674 4244 5686 4246
rect 5674 4236 5676 4244
rect 5684 4236 5686 4244
rect 5674 4184 5686 4236
rect 5674 4176 5676 4184
rect 5684 4176 5686 4184
rect 5674 4174 5686 4176
rect 5674 4144 5686 4146
rect 5674 4136 5676 4144
rect 5684 4136 5686 4144
rect 5578 3924 5590 3926
rect 5578 3916 5580 3924
rect 5588 3916 5590 3924
rect 5546 3764 5558 3766
rect 5546 3756 5548 3764
rect 5556 3756 5558 3764
rect 5546 3384 5558 3756
rect 5578 3624 5590 3916
rect 5674 3784 5686 4136
rect 5674 3776 5676 3784
rect 5684 3776 5686 3784
rect 5674 3774 5686 3776
rect 5706 4124 5718 4126
rect 5706 4116 5708 4124
rect 5716 4116 5718 4124
rect 5706 3864 5718 4116
rect 5834 4124 5846 4576
rect 6154 4564 6166 4566
rect 6154 4556 6156 4564
rect 6164 4556 6166 4564
rect 5994 4544 6006 4546
rect 5994 4536 5996 4544
rect 6004 4536 6006 4544
rect 5962 4504 5974 4506
rect 5962 4496 5964 4504
rect 5972 4496 5974 4504
rect 5898 4304 5910 4306
rect 5898 4296 5900 4304
rect 5908 4296 5910 4304
rect 5834 4116 5836 4124
rect 5844 4116 5846 4124
rect 5834 4114 5846 4116
rect 5866 4224 5878 4226
rect 5866 4216 5868 4224
rect 5876 4216 5878 4224
rect 5738 4104 5750 4106
rect 5738 4096 5740 4104
rect 5748 4096 5750 4104
rect 5738 3904 5750 4096
rect 5866 4084 5878 4216
rect 5866 4076 5868 4084
rect 5876 4076 5878 4084
rect 5866 4074 5878 4076
rect 5834 4064 5846 4066
rect 5834 4056 5836 4064
rect 5844 4056 5846 4064
rect 5738 3896 5740 3904
rect 5748 3896 5750 3904
rect 5738 3894 5750 3896
rect 5770 3904 5782 3906
rect 5770 3896 5772 3904
rect 5780 3896 5782 3904
rect 5706 3856 5708 3864
rect 5716 3856 5718 3864
rect 5642 3744 5654 3746
rect 5642 3736 5644 3744
rect 5652 3736 5654 3744
rect 5578 3616 5580 3624
rect 5588 3616 5590 3624
rect 5578 3614 5590 3616
rect 5610 3684 5622 3686
rect 5610 3676 5612 3684
rect 5620 3676 5622 3684
rect 5610 3484 5622 3676
rect 5610 3476 5612 3484
rect 5620 3476 5622 3484
rect 5546 3376 5548 3384
rect 5556 3376 5558 3384
rect 5546 3374 5558 3376
rect 5578 3404 5590 3406
rect 5578 3396 5580 3404
rect 5588 3396 5590 3404
rect 5514 3316 5516 3324
rect 5524 3316 5526 3324
rect 5514 3314 5526 3316
rect 5578 3244 5590 3396
rect 5578 3236 5580 3244
rect 5588 3236 5590 3244
rect 5578 3234 5590 3236
rect 5482 3056 5484 3064
rect 5492 3056 5494 3064
rect 5482 3054 5494 3056
rect 5546 3144 5558 3146
rect 5546 3136 5548 3144
rect 5556 3136 5558 3144
rect 5386 3016 5388 3024
rect 5396 3016 5398 3024
rect 5386 3014 5398 3016
rect 5546 3024 5558 3136
rect 5546 3016 5548 3024
rect 5556 3016 5558 3024
rect 5546 3014 5558 3016
rect 5482 2964 5494 2966
rect 5482 2956 5484 2964
rect 5492 2956 5494 2964
rect 5482 2664 5494 2956
rect 5610 2924 5622 3476
rect 5610 2916 5612 2924
rect 5620 2916 5622 2924
rect 5610 2914 5622 2916
rect 5642 3344 5654 3736
rect 5706 3704 5718 3856
rect 5706 3696 5708 3704
rect 5716 3696 5718 3704
rect 5706 3484 5718 3696
rect 5706 3476 5708 3484
rect 5716 3476 5718 3484
rect 5642 3336 5644 3344
rect 5652 3336 5654 3344
rect 5642 3104 5654 3336
rect 5642 3096 5644 3104
rect 5652 3096 5654 3104
rect 5642 3064 5654 3096
rect 5674 3444 5686 3446
rect 5674 3436 5676 3444
rect 5684 3436 5686 3444
rect 5674 3084 5686 3436
rect 5674 3076 5676 3084
rect 5684 3076 5686 3084
rect 5674 3074 5686 3076
rect 5642 3056 5644 3064
rect 5652 3056 5654 3064
rect 5642 2944 5654 3056
rect 5642 2936 5644 2944
rect 5652 2936 5654 2944
rect 5482 2656 5484 2664
rect 5492 2656 5494 2664
rect 5482 2654 5494 2656
rect 5578 2724 5590 2726
rect 5578 2716 5580 2724
rect 5588 2716 5590 2724
rect 5578 2624 5590 2716
rect 5610 2724 5622 2726
rect 5610 2716 5612 2724
rect 5620 2716 5622 2724
rect 5610 2644 5622 2716
rect 5610 2636 5612 2644
rect 5620 2636 5622 2644
rect 5610 2634 5622 2636
rect 5578 2616 5580 2624
rect 5588 2616 5590 2624
rect 5578 2614 5590 2616
rect 5354 2536 5356 2544
rect 5364 2536 5366 2544
rect 5354 2534 5366 2536
rect 5578 2564 5590 2566
rect 5578 2556 5580 2564
rect 5588 2556 5590 2564
rect 5322 2336 5324 2344
rect 5332 2336 5334 2344
rect 5322 2334 5334 2336
rect 5418 2484 5430 2486
rect 5418 2476 5420 2484
rect 5428 2476 5430 2484
rect 5034 2196 5036 2204
rect 5044 2196 5046 2204
rect 5034 2194 5046 2196
rect 5066 2304 5078 2306
rect 5066 2296 5068 2304
rect 5076 2296 5078 2304
rect 4938 2116 4940 2124
rect 4948 2116 4950 2124
rect 4938 2114 4950 2116
rect 5034 2124 5046 2126
rect 5034 2116 5036 2124
rect 5044 2116 5046 2124
rect 5002 2104 5014 2106
rect 5002 2096 5004 2104
rect 5012 2096 5014 2104
rect 5002 2004 5014 2096
rect 5002 1996 5004 2004
rect 5012 1996 5014 2004
rect 5002 1994 5014 1996
rect 4874 1896 4876 1904
rect 4884 1896 4886 1904
rect 4874 1894 4886 1896
rect 4906 1924 4918 1926
rect 4906 1916 4908 1924
rect 4916 1916 4918 1924
rect 4842 1856 4844 1864
rect 4852 1856 4854 1864
rect 4842 1854 4854 1856
rect 4778 1836 4780 1844
rect 4788 1836 4790 1844
rect 4778 1834 4790 1836
rect 4842 1824 4854 1826
rect 4842 1816 4844 1824
rect 4852 1816 4854 1824
rect 4664 1606 4666 1614
rect 4674 1606 4678 1614
rect 4686 1606 4690 1614
rect 4698 1606 4702 1614
rect 4710 1606 4712 1614
rect 4554 1276 4556 1284
rect 4564 1276 4566 1284
rect 4554 1274 4566 1276
rect 4586 1284 4598 1286
rect 4586 1276 4588 1284
rect 4596 1276 4598 1284
rect 4490 1216 4492 1224
rect 4500 1216 4502 1224
rect 4490 1214 4502 1216
rect 4586 1224 4598 1276
rect 4586 1216 4588 1224
rect 4596 1216 4598 1224
rect 4586 1214 4598 1216
rect 4664 1214 4712 1606
rect 4746 1664 4758 1666
rect 4746 1656 4748 1664
rect 4756 1656 4758 1664
rect 4746 1484 4758 1656
rect 4746 1476 4748 1484
rect 4756 1476 4758 1484
rect 4746 1474 4758 1476
rect 4810 1504 4822 1506
rect 4810 1496 4812 1504
rect 4820 1496 4822 1504
rect 4664 1206 4666 1214
rect 4674 1206 4678 1214
rect 4686 1206 4690 1214
rect 4698 1206 4702 1214
rect 4710 1206 4712 1214
rect 4778 1284 4790 1286
rect 4778 1276 4780 1284
rect 4788 1276 4790 1284
rect 4426 1156 4428 1164
rect 4436 1156 4438 1164
rect 4426 1154 4438 1156
rect 4554 1204 4566 1206
rect 4554 1196 4556 1204
rect 4564 1196 4566 1204
rect 4554 1144 4566 1196
rect 4554 1136 4556 1144
rect 4564 1136 4566 1144
rect 4554 1134 4566 1136
rect 4426 1124 4438 1126
rect 4426 1116 4428 1124
rect 4436 1116 4438 1124
rect 4426 1006 4438 1116
rect 4458 1124 4470 1126
rect 4458 1116 4460 1124
rect 4468 1116 4470 1124
rect 4458 1044 4470 1116
rect 4458 1036 4460 1044
rect 4468 1036 4470 1044
rect 4458 1034 4470 1036
rect 4522 1124 4534 1126
rect 4522 1116 4524 1124
rect 4532 1116 4534 1124
rect 4426 994 4502 1006
rect 4426 964 4438 966
rect 4426 956 4428 964
rect 4436 956 4438 964
rect 4426 884 4438 956
rect 4426 876 4428 884
rect 4436 876 4438 884
rect 4426 874 4438 876
rect 4458 964 4470 966
rect 4458 956 4460 964
rect 4468 956 4470 964
rect 4458 924 4470 956
rect 4458 916 4460 924
rect 4468 916 4470 924
rect 4394 796 4396 804
rect 4404 796 4406 804
rect 4394 794 4406 796
rect 4426 824 4438 826
rect 4426 816 4428 824
rect 4436 816 4438 824
rect 4426 624 4438 816
rect 4426 616 4428 624
rect 4436 616 4438 624
rect 4426 614 4438 616
rect 4458 624 4470 916
rect 4490 784 4502 994
rect 4490 776 4492 784
rect 4500 776 4502 784
rect 4490 774 4502 776
rect 4458 616 4460 624
rect 4468 616 4470 624
rect 4458 614 4470 616
rect 4362 436 4364 444
rect 4372 436 4374 444
rect 4362 434 4374 436
rect 4426 584 4438 586
rect 4426 576 4428 584
rect 4436 576 4438 584
rect 4426 484 4438 576
rect 4458 584 4470 586
rect 4458 576 4460 584
rect 4468 576 4470 584
rect 4458 566 4470 576
rect 4522 584 4534 1116
rect 4618 1124 4630 1126
rect 4618 1116 4620 1124
rect 4628 1116 4630 1124
rect 4554 1104 4566 1106
rect 4554 1096 4556 1104
rect 4564 1096 4566 1104
rect 4554 1024 4566 1096
rect 4554 1016 4556 1024
rect 4564 1016 4566 1024
rect 4554 1014 4566 1016
rect 4586 1084 4598 1086
rect 4586 1076 4588 1084
rect 4596 1076 4598 1084
rect 4586 904 4598 1076
rect 4618 984 4630 1116
rect 4618 976 4620 984
rect 4628 976 4630 984
rect 4618 974 4630 976
rect 4586 896 4588 904
rect 4596 896 4598 904
rect 4586 894 4598 896
rect 4618 924 4630 926
rect 4618 916 4620 924
rect 4628 916 4630 924
rect 4522 576 4524 584
rect 4532 576 4534 584
rect 4522 574 4534 576
rect 4554 884 4566 886
rect 4554 876 4556 884
rect 4564 876 4566 884
rect 4458 554 4502 566
rect 4426 476 4428 484
rect 4436 476 4438 484
rect 4394 424 4406 426
rect 4394 416 4396 424
rect 4404 416 4406 424
rect 4394 326 4406 416
rect 4330 156 4332 164
rect 4340 156 4342 164
rect 4330 154 4342 156
rect 4362 314 4406 326
rect 4298 136 4300 144
rect 4308 136 4310 144
rect 4298 134 4310 136
rect 4362 64 4374 314
rect 4394 284 4406 286
rect 4394 276 4396 284
rect 4404 276 4406 284
rect 4394 124 4406 276
rect 4394 116 4396 124
rect 4404 116 4406 124
rect 4394 114 4406 116
rect 4362 56 4364 64
rect 4372 56 4374 64
rect 4362 54 4374 56
rect 4426 64 4438 476
rect 4458 524 4470 526
rect 4458 516 4460 524
rect 4468 516 4470 524
rect 4458 486 4470 516
rect 4490 524 4502 554
rect 4490 516 4492 524
rect 4500 516 4502 524
rect 4490 514 4502 516
rect 4554 504 4566 876
rect 4586 824 4598 826
rect 4586 816 4588 824
rect 4596 816 4598 824
rect 4586 684 4598 816
rect 4586 676 4588 684
rect 4596 676 4598 684
rect 4586 674 4598 676
rect 4554 496 4556 504
rect 4564 496 4566 504
rect 4554 494 4566 496
rect 4618 624 4630 916
rect 4618 616 4620 624
rect 4628 616 4630 624
rect 4458 474 4534 486
rect 4490 404 4502 406
rect 4490 396 4492 404
rect 4500 396 4502 404
rect 4490 244 4502 396
rect 4522 404 4534 474
rect 4522 396 4524 404
rect 4532 396 4534 404
rect 4522 394 4534 396
rect 4554 404 4566 406
rect 4554 396 4556 404
rect 4564 396 4566 404
rect 4490 236 4492 244
rect 4500 236 4502 244
rect 4490 234 4502 236
rect 4522 324 4534 326
rect 4522 316 4524 324
rect 4532 316 4534 324
rect 4522 204 4534 316
rect 4554 324 4566 396
rect 4554 316 4556 324
rect 4564 316 4566 324
rect 4554 314 4566 316
rect 4586 324 4598 326
rect 4586 316 4588 324
rect 4596 316 4598 324
rect 4522 196 4524 204
rect 4532 196 4534 204
rect 4522 194 4534 196
rect 4554 284 4566 286
rect 4554 276 4556 284
rect 4564 276 4566 284
rect 4458 164 4502 166
rect 4458 156 4460 164
rect 4468 156 4502 164
rect 4458 154 4502 156
rect 4490 86 4502 154
rect 4490 84 4518 86
rect 4490 76 4508 84
rect 4516 76 4518 84
rect 4490 74 4518 76
rect 4426 56 4428 64
rect 4436 56 4438 64
rect 4426 54 4438 56
rect 4554 64 4566 276
rect 4586 264 4598 316
rect 4618 324 4630 616
rect 4618 316 4620 324
rect 4628 316 4630 324
rect 4618 314 4630 316
rect 4664 814 4712 1206
rect 4746 1204 4758 1206
rect 4746 1196 4748 1204
rect 4756 1196 4758 1204
rect 4746 1124 4758 1196
rect 4746 1116 4748 1124
rect 4756 1116 4758 1124
rect 4746 1114 4758 1116
rect 4778 1084 4790 1276
rect 4778 1076 4780 1084
rect 4788 1076 4790 1084
rect 4778 1074 4790 1076
rect 4664 806 4666 814
rect 4674 806 4678 814
rect 4686 806 4690 814
rect 4698 806 4702 814
rect 4710 806 4712 814
rect 4778 1004 4790 1006
rect 4778 996 4780 1004
rect 4788 996 4790 1004
rect 4664 414 4712 806
rect 4746 804 4758 806
rect 4746 796 4748 804
rect 4756 796 4758 804
rect 4746 724 4758 796
rect 4746 716 4748 724
rect 4756 716 4758 724
rect 4746 714 4758 716
rect 4746 684 4758 686
rect 4746 676 4748 684
rect 4756 676 4758 684
rect 4746 568 4758 676
rect 4778 644 4790 996
rect 4810 984 4822 1496
rect 4842 1404 4854 1816
rect 4906 1824 4918 1916
rect 4906 1816 4908 1824
rect 4916 1816 4918 1824
rect 4906 1814 4918 1816
rect 4970 1794 5014 1806
rect 4874 1784 4886 1786
rect 4874 1776 4876 1784
rect 4884 1776 4886 1784
rect 4874 1664 4886 1776
rect 4970 1744 4982 1794
rect 5002 1784 5014 1794
rect 5002 1776 5004 1784
rect 5012 1776 5014 1784
rect 5002 1774 5014 1776
rect 4970 1736 4972 1744
rect 4980 1736 4982 1744
rect 4970 1734 4982 1736
rect 4874 1656 4876 1664
rect 4884 1656 4886 1664
rect 4874 1654 4886 1656
rect 5034 1644 5046 2116
rect 5066 1924 5078 2296
rect 5130 2184 5142 2186
rect 5130 2176 5132 2184
rect 5140 2176 5142 2184
rect 5130 2104 5142 2176
rect 5130 2096 5132 2104
rect 5140 2096 5142 2104
rect 5130 2094 5142 2096
rect 5418 1984 5430 2476
rect 5418 1976 5420 1984
rect 5428 1976 5430 1984
rect 5418 1974 5430 1976
rect 5354 1944 5366 1946
rect 5354 1936 5356 1944
rect 5364 1936 5366 1944
rect 5354 1926 5366 1936
rect 5066 1916 5068 1924
rect 5076 1916 5078 1924
rect 5066 1914 5078 1916
rect 5098 1924 5110 1926
rect 5098 1916 5100 1924
rect 5108 1916 5110 1924
rect 5098 1864 5110 1916
rect 5322 1914 5366 1926
rect 5546 1924 5558 1926
rect 5546 1916 5548 1924
rect 5556 1916 5558 1924
rect 5098 1856 5100 1864
rect 5108 1856 5110 1864
rect 5098 1854 5110 1856
rect 5290 1904 5302 1906
rect 5290 1896 5292 1904
rect 5300 1896 5302 1904
rect 5034 1636 5036 1644
rect 5044 1636 5046 1644
rect 5034 1634 5046 1636
rect 5162 1564 5174 1566
rect 5162 1556 5164 1564
rect 5172 1556 5174 1564
rect 4938 1504 4950 1506
rect 4938 1496 4940 1504
rect 4948 1496 4950 1504
rect 4842 1396 4844 1404
rect 4852 1396 4854 1404
rect 4842 1394 4854 1396
rect 4874 1444 4886 1446
rect 4874 1436 4876 1444
rect 4884 1436 4886 1444
rect 4874 1284 4886 1436
rect 4874 1276 4876 1284
rect 4884 1276 4886 1284
rect 4874 1274 4886 1276
rect 4906 1284 4918 1286
rect 4906 1276 4908 1284
rect 4916 1276 4918 1284
rect 4842 1124 4854 1126
rect 4842 1116 4844 1124
rect 4852 1116 4854 1124
rect 4842 1064 4854 1116
rect 4842 1056 4844 1064
rect 4852 1056 4854 1064
rect 4842 1054 4854 1056
rect 4874 1064 4886 1066
rect 4874 1056 4876 1064
rect 4884 1056 4886 1064
rect 4810 976 4812 984
rect 4820 976 4822 984
rect 4810 974 4822 976
rect 4842 1004 4854 1006
rect 4842 996 4844 1004
rect 4852 996 4854 1004
rect 4778 636 4780 644
rect 4788 636 4790 644
rect 4778 634 4790 636
rect 4810 904 4822 906
rect 4810 896 4812 904
rect 4820 896 4822 904
rect 4810 684 4822 896
rect 4810 676 4812 684
rect 4820 676 4822 684
rect 4810 584 4822 676
rect 4810 576 4812 584
rect 4820 576 4822 584
rect 4810 574 4822 576
rect 4746 560 4748 568
rect 4756 560 4758 568
rect 4746 554 4758 560
rect 4746 540 4758 546
rect 4746 532 4748 540
rect 4756 532 4758 540
rect 4746 504 4758 532
rect 4746 496 4748 504
rect 4756 496 4758 504
rect 4746 494 4758 496
rect 4810 544 4822 546
rect 4810 536 4812 544
rect 4820 536 4822 544
rect 4664 406 4666 414
rect 4674 406 4678 414
rect 4686 406 4690 414
rect 4698 406 4702 414
rect 4710 406 4712 414
rect 4586 256 4588 264
rect 4596 256 4598 264
rect 4586 254 4598 256
rect 4554 56 4556 64
rect 4564 56 4566 64
rect 4554 54 4566 56
rect 4186 44 4214 46
rect 4186 36 4188 44
rect 4196 36 4214 44
rect 4186 34 4214 36
rect 4138 16 4140 24
rect 4148 16 4150 24
rect 4138 14 4150 16
rect 4664 14 4712 406
rect 4810 384 4822 536
rect 4810 376 4812 384
rect 4820 376 4822 384
rect 4810 374 4822 376
rect 4778 344 4790 346
rect 4778 336 4780 344
rect 4788 336 4790 344
rect 4778 304 4790 336
rect 4778 296 4780 304
rect 4788 296 4790 304
rect 4778 294 4790 296
rect 4842 264 4854 996
rect 4874 924 4886 1056
rect 4906 984 4918 1276
rect 4906 976 4908 984
rect 4916 976 4918 984
rect 4906 974 4918 976
rect 4874 916 4876 924
rect 4884 916 4886 924
rect 4874 914 4886 916
rect 4906 944 4918 946
rect 4906 936 4908 944
rect 4916 936 4918 944
rect 4874 644 4886 646
rect 4874 636 4876 644
rect 4884 636 4886 644
rect 4874 504 4886 636
rect 4906 524 4918 936
rect 4938 864 4950 1496
rect 5130 1464 5142 1466
rect 5130 1456 5132 1464
rect 5140 1456 5142 1464
rect 5034 1344 5046 1346
rect 5034 1336 5036 1344
rect 5044 1336 5046 1344
rect 5034 1326 5046 1336
rect 5002 1314 5046 1326
rect 5002 1304 5014 1314
rect 5002 1296 5004 1304
rect 5012 1296 5014 1304
rect 5002 1294 5014 1296
rect 5034 1264 5046 1266
rect 5034 1256 5036 1264
rect 5044 1256 5046 1264
rect 4970 1104 4982 1106
rect 4970 1096 4972 1104
rect 4980 1096 4982 1104
rect 4970 884 4982 1096
rect 5034 1004 5046 1256
rect 5098 1244 5110 1246
rect 5098 1236 5100 1244
rect 5108 1236 5110 1244
rect 5066 1084 5078 1086
rect 5066 1076 5068 1084
rect 5076 1076 5078 1084
rect 5066 1024 5078 1076
rect 5066 1016 5068 1024
rect 5076 1016 5078 1024
rect 5066 1014 5078 1016
rect 5034 996 5036 1004
rect 5044 996 5046 1004
rect 5034 994 5046 996
rect 5098 964 5110 1236
rect 5130 1124 5142 1456
rect 5162 1224 5174 1556
rect 5162 1216 5164 1224
rect 5172 1216 5174 1224
rect 5162 1214 5174 1216
rect 5194 1544 5206 1546
rect 5194 1536 5196 1544
rect 5204 1536 5206 1544
rect 5130 1116 5132 1124
rect 5140 1116 5142 1124
rect 5130 1114 5142 1116
rect 5162 1004 5174 1006
rect 5162 996 5164 1004
rect 5172 996 5174 1004
rect 5098 956 5100 964
rect 5108 956 5110 964
rect 5098 954 5110 956
rect 5130 964 5142 966
rect 5130 956 5132 964
rect 5140 956 5142 964
rect 5002 944 5014 946
rect 5002 936 5004 944
rect 5012 936 5014 944
rect 5002 904 5014 936
rect 5082 924 5110 926
rect 5082 916 5084 924
rect 5092 916 5110 924
rect 5082 914 5110 916
rect 5002 896 5004 904
rect 5012 896 5014 904
rect 5002 894 5014 896
rect 5066 904 5078 906
rect 5066 896 5068 904
rect 5076 896 5078 904
rect 4970 876 4972 884
rect 4980 876 4982 884
rect 4970 874 4982 876
rect 4938 856 4940 864
rect 4948 856 4950 864
rect 4938 854 4950 856
rect 5066 846 5078 896
rect 5098 884 5110 914
rect 5098 876 5100 884
rect 5108 876 5110 884
rect 5098 874 5110 876
rect 5050 844 5078 846
rect 5050 836 5052 844
rect 5060 836 5078 844
rect 5050 834 5078 836
rect 4970 804 4982 806
rect 4970 796 4972 804
rect 4980 796 4982 804
rect 4938 784 4950 786
rect 4938 776 4940 784
rect 4948 776 4950 784
rect 4938 584 4950 776
rect 4970 604 4982 796
rect 5066 784 5078 786
rect 5066 776 5068 784
rect 5076 776 5078 784
rect 5002 724 5014 726
rect 5002 716 5004 724
rect 5012 716 5014 724
rect 5002 624 5014 716
rect 5002 616 5004 624
rect 5012 616 5014 624
rect 5002 614 5014 616
rect 4970 596 4972 604
rect 4980 596 4982 604
rect 4970 594 4982 596
rect 5066 604 5078 776
rect 5066 596 5068 604
rect 5076 596 5078 604
rect 5066 594 5078 596
rect 5098 744 5110 746
rect 5098 736 5100 744
rect 5108 736 5110 744
rect 4938 576 4940 584
rect 4948 576 4950 584
rect 4938 574 4950 576
rect 5098 564 5110 736
rect 5098 556 5100 564
rect 5108 556 5110 564
rect 4906 516 4908 524
rect 4916 516 4918 524
rect 4906 514 4918 516
rect 5002 524 5014 526
rect 5002 516 5004 524
rect 5012 516 5014 524
rect 4874 496 4876 504
rect 4884 496 4886 504
rect 4874 494 4886 496
rect 4970 464 4982 466
rect 4970 456 4972 464
rect 4980 456 4982 464
rect 4970 424 4982 456
rect 4970 416 4972 424
rect 4980 416 4982 424
rect 4970 414 4982 416
rect 4842 256 4844 264
rect 4852 256 4854 264
rect 4842 254 4854 256
rect 4874 404 4886 406
rect 4874 396 4876 404
rect 4884 396 4886 404
rect 4810 244 4822 246
rect 4810 236 4812 244
rect 4820 236 4822 244
rect 4810 124 4822 236
rect 4874 164 4886 396
rect 5002 304 5014 516
rect 5066 524 5078 526
rect 5066 516 5068 524
rect 5076 516 5078 524
rect 5034 464 5046 466
rect 5034 456 5036 464
rect 5044 456 5046 464
rect 5034 404 5046 456
rect 5034 396 5036 404
rect 5044 396 5046 404
rect 5034 394 5046 396
rect 5002 296 5004 304
rect 5012 296 5014 304
rect 5002 294 5014 296
rect 4874 156 4876 164
rect 4884 156 4886 164
rect 4874 154 4886 156
rect 4938 264 4950 266
rect 4938 256 4940 264
rect 4948 256 4950 264
rect 4810 116 4812 124
rect 4820 116 4822 124
rect 4810 114 4822 116
rect 4938 86 4950 256
rect 5034 264 5046 266
rect 5034 256 5036 264
rect 5044 256 5046 264
rect 5034 184 5046 256
rect 5034 176 5036 184
rect 5044 176 5046 184
rect 5034 174 5046 176
rect 5002 164 5014 166
rect 5002 156 5004 164
rect 5012 156 5014 164
rect 4938 84 4966 86
rect 4938 76 4956 84
rect 4964 76 4966 84
rect 4938 74 4966 76
rect 5002 64 5014 156
rect 5002 56 5004 64
rect 5012 56 5014 64
rect 5002 54 5014 56
rect 5034 144 5046 146
rect 5034 136 5036 144
rect 5044 136 5046 144
rect 5034 64 5046 136
rect 5066 104 5078 516
rect 5098 304 5110 556
rect 5130 524 5142 956
rect 5162 924 5174 996
rect 5162 916 5164 924
rect 5172 916 5174 924
rect 5162 914 5174 916
rect 5194 704 5206 1536
rect 5258 1544 5270 1546
rect 5258 1536 5260 1544
rect 5268 1536 5270 1544
rect 5258 1484 5270 1536
rect 5258 1476 5260 1484
rect 5268 1476 5270 1484
rect 5258 1474 5270 1476
rect 5226 1324 5238 1326
rect 5226 1316 5228 1324
rect 5236 1316 5238 1324
rect 5226 1044 5238 1316
rect 5290 1284 5302 1896
rect 5322 1884 5334 1914
rect 5322 1876 5324 1884
rect 5332 1876 5334 1884
rect 5322 1874 5334 1876
rect 5450 1884 5462 1886
rect 5450 1876 5452 1884
rect 5460 1876 5462 1884
rect 5290 1276 5292 1284
rect 5300 1276 5302 1284
rect 5290 1274 5302 1276
rect 5322 1744 5334 1746
rect 5322 1736 5324 1744
rect 5332 1736 5334 1744
rect 5322 1484 5334 1736
rect 5450 1704 5462 1876
rect 5450 1696 5452 1704
rect 5460 1696 5462 1704
rect 5450 1664 5462 1696
rect 5450 1656 5452 1664
rect 5460 1656 5462 1664
rect 5450 1654 5462 1656
rect 5514 1784 5526 1786
rect 5514 1776 5516 1784
rect 5524 1776 5526 1784
rect 5482 1644 5494 1646
rect 5482 1636 5484 1644
rect 5492 1636 5494 1644
rect 5322 1476 5324 1484
rect 5332 1476 5334 1484
rect 5290 1244 5302 1246
rect 5290 1236 5292 1244
rect 5300 1236 5302 1244
rect 5226 1036 5228 1044
rect 5236 1036 5238 1044
rect 5226 1034 5238 1036
rect 5258 1164 5270 1166
rect 5258 1156 5260 1164
rect 5268 1156 5270 1164
rect 5226 964 5238 966
rect 5226 956 5228 964
rect 5236 956 5238 964
rect 5226 904 5238 956
rect 5226 896 5228 904
rect 5236 896 5238 904
rect 5226 894 5238 896
rect 5258 784 5270 1156
rect 5290 944 5302 1236
rect 5322 1084 5334 1476
rect 5386 1624 5398 1626
rect 5386 1616 5388 1624
rect 5396 1616 5398 1624
rect 5322 1076 5324 1084
rect 5332 1076 5334 1084
rect 5322 1074 5334 1076
rect 5354 1324 5366 1326
rect 5354 1316 5356 1324
rect 5364 1316 5366 1324
rect 5290 936 5292 944
rect 5300 936 5302 944
rect 5290 934 5302 936
rect 5322 964 5334 966
rect 5322 956 5324 964
rect 5332 956 5334 964
rect 5322 824 5334 956
rect 5354 864 5366 1316
rect 5386 1024 5398 1616
rect 5482 1584 5494 1636
rect 5482 1576 5484 1584
rect 5492 1576 5494 1584
rect 5482 1574 5494 1576
rect 5514 1504 5526 1776
rect 5514 1496 5516 1504
rect 5524 1496 5526 1504
rect 5514 1494 5526 1496
rect 5482 1444 5494 1446
rect 5482 1436 5484 1444
rect 5492 1436 5494 1444
rect 5450 1284 5462 1286
rect 5450 1276 5452 1284
rect 5460 1276 5462 1284
rect 5386 1016 5388 1024
rect 5396 1016 5398 1024
rect 5386 1014 5398 1016
rect 5418 1064 5430 1066
rect 5418 1056 5420 1064
rect 5428 1056 5430 1064
rect 5418 964 5430 1056
rect 5418 956 5420 964
rect 5428 956 5430 964
rect 5418 954 5430 956
rect 5354 856 5356 864
rect 5364 856 5366 864
rect 5354 854 5366 856
rect 5386 884 5398 886
rect 5386 876 5388 884
rect 5396 876 5398 884
rect 5386 864 5398 876
rect 5386 856 5388 864
rect 5396 856 5398 864
rect 5322 816 5324 824
rect 5332 816 5334 824
rect 5322 814 5334 816
rect 5258 776 5260 784
rect 5268 776 5270 784
rect 5258 774 5270 776
rect 5354 784 5366 786
rect 5354 776 5356 784
rect 5364 776 5366 784
rect 5194 696 5196 704
rect 5204 696 5206 704
rect 5194 694 5206 696
rect 5258 704 5270 706
rect 5258 696 5260 704
rect 5268 696 5270 704
rect 5226 664 5238 666
rect 5226 656 5228 664
rect 5236 656 5238 664
rect 5226 604 5238 656
rect 5226 596 5228 604
rect 5236 596 5238 604
rect 5226 594 5238 596
rect 5258 604 5270 696
rect 5354 704 5366 776
rect 5354 696 5356 704
rect 5364 696 5366 704
rect 5354 694 5366 696
rect 5306 684 5350 686
rect 5306 676 5308 684
rect 5316 676 5340 684
rect 5348 676 5350 684
rect 5306 674 5350 676
rect 5258 596 5260 604
rect 5268 596 5270 604
rect 5258 594 5270 596
rect 5290 664 5302 666
rect 5290 656 5292 664
rect 5300 656 5302 664
rect 5130 516 5132 524
rect 5140 516 5142 524
rect 5130 514 5142 516
rect 5162 584 5174 586
rect 5162 576 5164 584
rect 5172 576 5174 584
rect 5098 296 5100 304
rect 5108 296 5110 304
rect 5098 294 5110 296
rect 5130 304 5142 306
rect 5130 296 5132 304
rect 5140 296 5142 304
rect 5130 164 5142 296
rect 5162 284 5174 576
rect 5290 564 5302 656
rect 5290 556 5292 564
rect 5300 556 5302 564
rect 5290 554 5302 556
rect 5322 664 5334 666
rect 5322 656 5324 664
rect 5332 656 5334 664
rect 5226 544 5238 546
rect 5226 536 5228 544
rect 5236 536 5238 544
rect 5226 384 5238 536
rect 5226 376 5228 384
rect 5236 376 5238 384
rect 5226 374 5238 376
rect 5258 544 5270 546
rect 5258 536 5260 544
rect 5268 536 5270 544
rect 5162 276 5164 284
rect 5172 276 5174 284
rect 5162 274 5174 276
rect 5130 156 5132 164
rect 5140 156 5142 164
rect 5130 154 5142 156
rect 5194 164 5206 166
rect 5194 156 5196 164
rect 5204 156 5206 164
rect 5066 96 5068 104
rect 5076 96 5078 104
rect 5066 94 5078 96
rect 5194 84 5206 156
rect 5194 76 5196 84
rect 5204 76 5206 84
rect 5194 74 5206 76
rect 5034 56 5036 64
rect 5044 56 5046 64
rect 5034 54 5046 56
rect 5258 44 5270 536
rect 5322 464 5334 656
rect 5354 624 5366 626
rect 5354 616 5356 624
rect 5364 616 5366 624
rect 5354 504 5366 616
rect 5386 624 5398 856
rect 5386 616 5388 624
rect 5396 616 5398 624
rect 5386 614 5398 616
rect 5418 824 5430 826
rect 5418 816 5420 824
rect 5428 816 5430 824
rect 5418 624 5430 816
rect 5418 616 5420 624
rect 5428 616 5430 624
rect 5418 614 5430 616
rect 5450 524 5462 1276
rect 5482 1224 5494 1436
rect 5482 1216 5484 1224
rect 5492 1216 5494 1224
rect 5482 1214 5494 1216
rect 5514 1324 5526 1326
rect 5514 1316 5516 1324
rect 5524 1316 5526 1324
rect 5514 1084 5526 1316
rect 5546 1104 5558 1916
rect 5578 1504 5590 2556
rect 5642 2544 5654 2936
rect 5642 2536 5644 2544
rect 5652 2536 5654 2544
rect 5610 2044 5622 2046
rect 5610 2036 5612 2044
rect 5620 2036 5622 2044
rect 5610 1724 5622 2036
rect 5610 1716 5612 1724
rect 5620 1716 5622 1724
rect 5610 1714 5622 1716
rect 5578 1496 5580 1504
rect 5588 1496 5590 1504
rect 5578 1494 5590 1496
rect 5610 1664 5622 1666
rect 5610 1656 5612 1664
rect 5620 1656 5622 1664
rect 5546 1096 5548 1104
rect 5556 1096 5558 1104
rect 5546 1094 5558 1096
rect 5578 1464 5590 1466
rect 5578 1456 5580 1464
rect 5588 1456 5590 1464
rect 5514 1076 5516 1084
rect 5524 1076 5526 1084
rect 5514 1074 5526 1076
rect 5482 1064 5494 1066
rect 5482 1056 5484 1064
rect 5492 1056 5494 1064
rect 5482 948 5494 1056
rect 5482 940 5484 948
rect 5492 940 5494 948
rect 5482 934 5494 940
rect 5514 964 5526 966
rect 5514 956 5516 964
rect 5524 956 5526 964
rect 5482 920 5494 926
rect 5482 912 5484 920
rect 5492 912 5494 920
rect 5482 744 5494 912
rect 5482 736 5484 744
rect 5492 736 5494 744
rect 5482 734 5494 736
rect 5450 516 5452 524
rect 5460 516 5462 524
rect 5450 514 5462 516
rect 5482 704 5494 706
rect 5482 696 5484 704
rect 5492 696 5494 704
rect 5354 496 5356 504
rect 5364 496 5366 504
rect 5354 494 5366 496
rect 5322 456 5324 464
rect 5332 456 5334 464
rect 5322 454 5334 456
rect 5354 464 5366 466
rect 5354 456 5356 464
rect 5364 456 5366 464
rect 5354 424 5366 456
rect 5354 416 5356 424
rect 5364 416 5366 424
rect 5354 324 5366 416
rect 5354 316 5356 324
rect 5364 316 5366 324
rect 5354 314 5366 316
rect 5418 464 5430 466
rect 5418 456 5420 464
rect 5428 456 5430 464
rect 5418 264 5430 456
rect 5418 256 5420 264
rect 5428 256 5430 264
rect 5418 254 5430 256
rect 5450 264 5462 266
rect 5450 256 5452 264
rect 5460 256 5462 264
rect 5274 204 5302 206
rect 5274 196 5276 204
rect 5284 196 5302 204
rect 5274 194 5302 196
rect 5290 124 5302 194
rect 5418 204 5430 206
rect 5418 196 5420 204
rect 5428 196 5430 204
rect 5354 184 5366 186
rect 5354 176 5356 184
rect 5364 176 5366 184
rect 5290 116 5292 124
rect 5300 116 5302 124
rect 5290 114 5302 116
rect 5322 124 5334 126
rect 5322 116 5324 124
rect 5332 116 5334 124
rect 5322 86 5334 116
rect 5258 36 5260 44
rect 5268 36 5270 44
rect 5258 34 5270 36
rect 5290 74 5334 86
rect 5290 44 5302 74
rect 5290 36 5292 44
rect 5300 36 5302 44
rect 5290 34 5302 36
rect 5354 24 5366 176
rect 5354 16 5356 24
rect 5364 16 5366 24
rect 5354 14 5366 16
rect 5386 124 5398 126
rect 5386 116 5388 124
rect 5396 116 5398 124
rect 5386 24 5398 116
rect 5418 84 5430 196
rect 5418 76 5420 84
rect 5428 76 5430 84
rect 5418 74 5430 76
rect 5450 64 5462 256
rect 5450 56 5452 64
rect 5460 56 5462 64
rect 5450 54 5462 56
rect 5386 16 5388 24
rect 5396 16 5398 24
rect 5386 14 5398 16
rect 5482 24 5494 696
rect 5514 704 5526 956
rect 5514 696 5516 704
rect 5524 696 5526 704
rect 5514 694 5526 696
rect 5514 604 5526 606
rect 5514 596 5516 604
rect 5524 596 5526 604
rect 5514 484 5526 596
rect 5514 476 5516 484
rect 5524 476 5526 484
rect 5514 474 5526 476
rect 5546 564 5558 566
rect 5546 556 5548 564
rect 5556 556 5558 564
rect 5546 424 5558 556
rect 5546 416 5548 424
rect 5556 416 5558 424
rect 5546 414 5558 416
rect 5578 144 5590 1456
rect 5610 1324 5622 1656
rect 5610 1316 5612 1324
rect 5620 1316 5622 1324
rect 5610 1314 5622 1316
rect 5610 1224 5622 1226
rect 5610 1216 5612 1224
rect 5620 1216 5622 1224
rect 5610 1024 5622 1216
rect 5610 1016 5612 1024
rect 5620 1016 5622 1024
rect 5610 1014 5622 1016
rect 5610 964 5622 966
rect 5610 956 5612 964
rect 5620 956 5622 964
rect 5610 484 5622 956
rect 5610 476 5612 484
rect 5620 476 5622 484
rect 5610 474 5622 476
rect 5642 184 5654 2536
rect 5674 2784 5686 2786
rect 5674 2776 5676 2784
rect 5684 2776 5686 2784
rect 5674 2344 5686 2776
rect 5674 2336 5676 2344
rect 5684 2336 5686 2344
rect 5674 2334 5686 2336
rect 5706 2724 5718 3476
rect 5738 3724 5750 3726
rect 5738 3716 5740 3724
rect 5748 3716 5750 3724
rect 5738 3464 5750 3716
rect 5770 3544 5782 3896
rect 5834 3824 5846 4056
rect 5834 3816 5836 3824
rect 5844 3816 5846 3824
rect 5834 3814 5846 3816
rect 5770 3536 5772 3544
rect 5780 3536 5782 3544
rect 5770 3534 5782 3536
rect 5802 3784 5814 3786
rect 5802 3776 5804 3784
rect 5812 3776 5814 3784
rect 5802 3524 5814 3776
rect 5834 3784 5846 3786
rect 5834 3776 5836 3784
rect 5844 3776 5846 3784
rect 5834 3704 5846 3776
rect 5834 3696 5836 3704
rect 5844 3696 5846 3704
rect 5834 3694 5846 3696
rect 5898 3764 5910 4296
rect 5930 4264 5942 4266
rect 5930 4256 5932 4264
rect 5940 4256 5942 4264
rect 5930 4164 5942 4256
rect 5930 4156 5932 4164
rect 5940 4156 5942 4164
rect 5930 3944 5942 4156
rect 5930 3936 5932 3944
rect 5940 3936 5942 3944
rect 5930 3934 5942 3936
rect 5898 3756 5900 3764
rect 5908 3756 5910 3764
rect 5802 3516 5804 3524
rect 5812 3516 5814 3524
rect 5802 3514 5814 3516
rect 5834 3624 5846 3626
rect 5834 3616 5836 3624
rect 5844 3616 5846 3624
rect 5834 3524 5846 3616
rect 5834 3516 5836 3524
rect 5844 3516 5846 3524
rect 5834 3514 5846 3516
rect 5866 3544 5878 3546
rect 5866 3536 5868 3544
rect 5876 3536 5878 3544
rect 5738 3456 5740 3464
rect 5748 3456 5750 3464
rect 5738 3454 5750 3456
rect 5834 3424 5846 3426
rect 5834 3416 5836 3424
rect 5844 3416 5846 3424
rect 5738 3404 5750 3406
rect 5738 3396 5740 3404
rect 5748 3396 5750 3404
rect 5738 2924 5750 3396
rect 5802 3184 5814 3186
rect 5802 3176 5804 3184
rect 5812 3176 5814 3184
rect 5802 2984 5814 3176
rect 5802 2976 5804 2984
rect 5812 2976 5814 2984
rect 5802 2974 5814 2976
rect 5738 2916 5740 2924
rect 5748 2916 5750 2924
rect 5738 2744 5750 2916
rect 5802 2944 5814 2946
rect 5802 2936 5804 2944
rect 5812 2936 5814 2944
rect 5802 2884 5814 2936
rect 5802 2876 5804 2884
rect 5812 2876 5814 2884
rect 5802 2874 5814 2876
rect 5738 2736 5740 2744
rect 5748 2736 5750 2744
rect 5738 2734 5750 2736
rect 5770 2844 5782 2846
rect 5770 2836 5772 2844
rect 5780 2836 5782 2844
rect 5706 2716 5708 2724
rect 5716 2716 5718 2724
rect 5706 2704 5718 2716
rect 5706 2696 5708 2704
rect 5716 2696 5718 2704
rect 5674 2304 5686 2306
rect 5674 2296 5676 2304
rect 5684 2296 5686 2304
rect 5674 2224 5686 2296
rect 5674 2216 5676 2224
rect 5684 2216 5686 2224
rect 5674 1004 5686 2216
rect 5706 1904 5718 2696
rect 5706 1896 5708 1904
rect 5716 1896 5718 1904
rect 5706 1894 5718 1896
rect 5738 2664 5750 2666
rect 5738 2656 5740 2664
rect 5748 2656 5750 2664
rect 5738 1944 5750 2656
rect 5770 2564 5782 2836
rect 5802 2824 5814 2826
rect 5802 2816 5804 2824
rect 5812 2816 5814 2824
rect 5802 2624 5814 2816
rect 5802 2616 5804 2624
rect 5812 2616 5814 2624
rect 5802 2614 5814 2616
rect 5770 2556 5772 2564
rect 5780 2556 5782 2564
rect 5770 2554 5782 2556
rect 5770 2514 5814 2526
rect 5834 2524 5846 3416
rect 5834 2516 5836 2524
rect 5844 2516 5846 2524
rect 5834 2514 5846 2516
rect 5770 2484 5782 2514
rect 5802 2504 5814 2514
rect 5802 2496 5804 2504
rect 5812 2496 5814 2504
rect 5802 2494 5814 2496
rect 5770 2476 5772 2484
rect 5780 2476 5782 2484
rect 5770 2474 5782 2476
rect 5802 2404 5814 2406
rect 5802 2396 5804 2404
rect 5812 2396 5814 2404
rect 5738 1936 5740 1944
rect 5748 1936 5750 1944
rect 5706 1864 5718 1866
rect 5706 1856 5708 1864
rect 5716 1856 5718 1864
rect 5706 1684 5718 1856
rect 5706 1676 5708 1684
rect 5716 1676 5718 1684
rect 5706 1674 5718 1676
rect 5674 996 5676 1004
rect 5684 996 5686 1004
rect 5674 994 5686 996
rect 5706 1504 5718 1506
rect 5706 1496 5708 1504
rect 5716 1496 5718 1504
rect 5674 864 5686 866
rect 5674 856 5676 864
rect 5684 856 5686 864
rect 5674 344 5686 856
rect 5674 336 5676 344
rect 5684 336 5686 344
rect 5674 334 5686 336
rect 5642 176 5644 184
rect 5652 176 5654 184
rect 5642 174 5654 176
rect 5674 284 5686 286
rect 5674 276 5676 284
rect 5684 276 5686 284
rect 5578 136 5580 144
rect 5588 136 5590 144
rect 5578 134 5590 136
rect 5674 104 5686 276
rect 5706 124 5718 1496
rect 5706 116 5708 124
rect 5716 116 5718 124
rect 5706 114 5718 116
rect 5738 124 5750 1936
rect 5770 2344 5782 2346
rect 5770 2336 5772 2344
rect 5780 2336 5782 2344
rect 5770 1564 5782 2336
rect 5802 2264 5814 2396
rect 5802 2256 5804 2264
rect 5812 2256 5814 2264
rect 5802 2254 5814 2256
rect 5834 2284 5846 2286
rect 5834 2276 5836 2284
rect 5844 2276 5846 2284
rect 5770 1556 5772 1564
rect 5780 1556 5782 1564
rect 5770 1554 5782 1556
rect 5802 2184 5814 2186
rect 5802 2176 5804 2184
rect 5812 2176 5814 2184
rect 5770 1524 5782 1526
rect 5770 1516 5772 1524
rect 5780 1516 5782 1524
rect 5770 1404 5782 1516
rect 5770 1396 5772 1404
rect 5780 1396 5782 1404
rect 5770 1394 5782 1396
rect 5770 1204 5782 1206
rect 5770 1196 5772 1204
rect 5780 1196 5782 1204
rect 5770 868 5782 1196
rect 5770 860 5772 868
rect 5780 860 5782 868
rect 5770 854 5782 860
rect 5770 840 5782 846
rect 5770 832 5772 840
rect 5780 832 5782 840
rect 5770 424 5782 832
rect 5770 416 5772 424
rect 5780 416 5782 424
rect 5770 414 5782 416
rect 5770 364 5782 366
rect 5770 356 5772 364
rect 5780 356 5782 364
rect 5770 284 5782 356
rect 5770 276 5772 284
rect 5780 276 5782 284
rect 5770 274 5782 276
rect 5802 164 5814 2176
rect 5834 2184 5846 2276
rect 5834 2176 5836 2184
rect 5844 2176 5846 2184
rect 5834 2174 5846 2176
rect 5834 1744 5846 1746
rect 5834 1736 5836 1744
rect 5844 1736 5846 1744
rect 5834 1464 5846 1736
rect 5834 1456 5836 1464
rect 5844 1456 5846 1464
rect 5834 1454 5846 1456
rect 5834 1364 5846 1366
rect 5834 1356 5836 1364
rect 5844 1356 5846 1364
rect 5834 1164 5846 1356
rect 5834 1156 5836 1164
rect 5844 1156 5846 1164
rect 5834 1154 5846 1156
rect 5834 1124 5846 1126
rect 5834 1116 5836 1124
rect 5844 1116 5846 1124
rect 5834 1024 5846 1116
rect 5866 1104 5878 3536
rect 5866 1096 5868 1104
rect 5876 1096 5878 1104
rect 5866 1094 5878 1096
rect 5898 3324 5910 3756
rect 5930 3764 5942 3766
rect 5930 3756 5932 3764
rect 5940 3756 5942 3764
rect 5930 3504 5942 3756
rect 5962 3544 5974 4496
rect 5962 3536 5964 3544
rect 5972 3536 5974 3544
rect 5962 3534 5974 3536
rect 5930 3496 5932 3504
rect 5940 3496 5942 3504
rect 5930 3494 5942 3496
rect 5962 3484 5974 3486
rect 5962 3476 5964 3484
rect 5972 3476 5974 3484
rect 5962 3444 5974 3476
rect 5962 3436 5964 3444
rect 5972 3436 5974 3444
rect 5962 3434 5974 3436
rect 5898 3316 5900 3324
rect 5908 3316 5910 3324
rect 5898 3084 5910 3316
rect 5962 3404 5974 3406
rect 5962 3396 5964 3404
rect 5972 3396 5974 3404
rect 5930 3164 5942 3166
rect 5930 3156 5932 3164
rect 5940 3156 5942 3164
rect 5930 3104 5942 3156
rect 5930 3096 5932 3104
rect 5940 3096 5942 3104
rect 5930 3094 5942 3096
rect 5898 3076 5900 3084
rect 5908 3076 5910 3084
rect 5898 2704 5910 3076
rect 5898 2696 5900 2704
rect 5908 2696 5910 2704
rect 5834 1016 5836 1024
rect 5844 1016 5846 1024
rect 5834 1014 5846 1016
rect 5866 1024 5878 1026
rect 5866 1016 5868 1024
rect 5876 1016 5878 1024
rect 5834 984 5846 986
rect 5834 976 5836 984
rect 5844 976 5846 984
rect 5834 544 5846 976
rect 5834 536 5836 544
rect 5844 536 5846 544
rect 5834 534 5846 536
rect 5866 504 5878 1016
rect 5898 924 5910 2696
rect 5930 2764 5942 2766
rect 5930 2756 5932 2764
rect 5940 2756 5942 2764
rect 5930 2664 5942 2756
rect 5930 2656 5932 2664
rect 5940 2656 5942 2664
rect 5930 2654 5942 2656
rect 5930 2604 5942 2606
rect 5930 2596 5932 2604
rect 5940 2596 5942 2604
rect 5930 2284 5942 2596
rect 5930 2276 5932 2284
rect 5940 2276 5942 2284
rect 5930 2274 5942 2276
rect 5930 1864 5942 1866
rect 5930 1856 5932 1864
rect 5940 1856 5942 1864
rect 5930 1444 5942 1856
rect 5930 1436 5932 1444
rect 5940 1436 5942 1444
rect 5930 1434 5942 1436
rect 5930 1404 5942 1406
rect 5930 1396 5932 1404
rect 5940 1396 5942 1404
rect 5930 944 5942 1396
rect 5962 1404 5974 3396
rect 5962 1396 5964 1404
rect 5972 1396 5974 1404
rect 5962 1394 5974 1396
rect 5994 1484 6006 4536
rect 6154 4504 6166 4556
rect 6154 4496 6156 4504
rect 6164 4496 6166 4504
rect 6154 4494 6166 4496
rect 6154 4464 6166 4466
rect 6154 4456 6156 4464
rect 6164 4456 6166 4464
rect 6026 4264 6038 4266
rect 6026 4256 6028 4264
rect 6036 4256 6038 4264
rect 6026 4084 6038 4256
rect 6122 4264 6134 4266
rect 6122 4256 6124 4264
rect 6132 4256 6134 4264
rect 6122 4164 6134 4256
rect 6122 4156 6124 4164
rect 6132 4156 6134 4164
rect 6026 4076 6028 4084
rect 6036 4076 6038 4084
rect 6026 3844 6038 4076
rect 6090 4084 6102 4086
rect 6090 4076 6092 4084
rect 6100 4076 6102 4084
rect 6026 3836 6028 3844
rect 6036 3836 6038 3844
rect 6026 3834 6038 3836
rect 6058 3984 6070 3986
rect 6058 3976 6060 3984
rect 6068 3976 6070 3984
rect 6058 3784 6070 3976
rect 6058 3776 6060 3784
rect 6068 3776 6070 3784
rect 6058 3774 6070 3776
rect 6026 3704 6038 3706
rect 6026 3696 6028 3704
rect 6036 3696 6038 3704
rect 6026 2584 6038 3696
rect 6090 3604 6102 4076
rect 6122 4044 6134 4156
rect 6122 4036 6124 4044
rect 6132 4036 6134 4044
rect 6122 4034 6134 4036
rect 6154 3924 6166 4456
rect 6250 4344 6262 4346
rect 6250 4336 6252 4344
rect 6260 4336 6262 4344
rect 6154 3916 6156 3924
rect 6164 3916 6166 3924
rect 6154 3914 6166 3916
rect 6186 4164 6198 4166
rect 6186 4156 6188 4164
rect 6196 4156 6198 4164
rect 6122 3904 6134 3906
rect 6122 3896 6124 3904
rect 6132 3896 6134 3904
rect 6122 3784 6134 3896
rect 6186 3884 6198 4156
rect 6186 3876 6188 3884
rect 6196 3876 6198 3884
rect 6186 3874 6198 3876
rect 6218 4124 6230 4126
rect 6218 4116 6220 4124
rect 6228 4116 6230 4124
rect 6122 3776 6124 3784
rect 6132 3776 6134 3784
rect 6122 3774 6134 3776
rect 6154 3824 6166 3826
rect 6154 3816 6156 3824
rect 6164 3816 6166 3824
rect 6154 3724 6166 3816
rect 6154 3716 6156 3724
rect 6164 3716 6166 3724
rect 6154 3714 6166 3716
rect 6186 3804 6198 3806
rect 6186 3796 6188 3804
rect 6196 3796 6198 3804
rect 6090 3596 6092 3604
rect 6100 3596 6102 3604
rect 6090 3594 6102 3596
rect 6122 3684 6134 3686
rect 6122 3676 6124 3684
rect 6132 3676 6134 3684
rect 6122 3464 6134 3676
rect 6122 3456 6124 3464
rect 6132 3456 6134 3464
rect 6122 3454 6134 3456
rect 6026 2576 6028 2584
rect 6036 2576 6038 2584
rect 6026 2574 6038 2576
rect 6090 3444 6102 3446
rect 6090 3436 6092 3444
rect 6100 3436 6102 3444
rect 6090 2664 6102 3436
rect 6186 3384 6198 3796
rect 6186 3376 6188 3384
rect 6196 3376 6198 3384
rect 6186 3374 6198 3376
rect 6122 3364 6134 3366
rect 6122 3356 6124 3364
rect 6132 3356 6134 3364
rect 6122 3284 6134 3356
rect 6186 3344 6198 3346
rect 6186 3336 6188 3344
rect 6196 3336 6198 3344
rect 6122 3276 6124 3284
rect 6132 3276 6134 3284
rect 6122 3274 6134 3276
rect 6154 3304 6166 3306
rect 6154 3296 6156 3304
rect 6164 3296 6166 3304
rect 6122 3024 6134 3026
rect 6122 3016 6124 3024
rect 6132 3016 6134 3024
rect 6122 2724 6134 3016
rect 6154 2744 6166 3296
rect 6186 3304 6198 3336
rect 6186 3296 6188 3304
rect 6196 3296 6198 3304
rect 6186 3294 6198 3296
rect 6186 3124 6198 3126
rect 6186 3116 6188 3124
rect 6196 3116 6198 3124
rect 6186 2964 6198 3116
rect 6186 2956 6188 2964
rect 6196 2956 6198 2964
rect 6186 2904 6198 2956
rect 6186 2896 6188 2904
rect 6196 2896 6198 2904
rect 6186 2894 6198 2896
rect 6154 2736 6156 2744
rect 6164 2736 6166 2744
rect 6154 2734 6166 2736
rect 6122 2716 6124 2724
rect 6132 2716 6134 2724
rect 6122 2714 6134 2716
rect 6090 2656 6092 2664
rect 6100 2656 6102 2664
rect 6058 2524 6070 2526
rect 6058 2516 6060 2524
rect 6068 2516 6070 2524
rect 6026 2444 6038 2446
rect 6026 2436 6028 2444
rect 6036 2436 6038 2444
rect 6026 2144 6038 2436
rect 6058 2344 6070 2516
rect 6058 2336 6060 2344
rect 6068 2336 6070 2344
rect 6058 2334 6070 2336
rect 6026 2136 6028 2144
rect 6036 2136 6038 2144
rect 6026 2134 6038 2136
rect 5994 1476 5996 1484
rect 6004 1476 6006 1484
rect 5962 1344 5974 1346
rect 5962 1336 5964 1344
rect 5972 1336 5974 1344
rect 5962 1144 5974 1336
rect 5962 1136 5964 1144
rect 5972 1136 5974 1144
rect 5962 1134 5974 1136
rect 5994 1344 6006 1476
rect 6026 2084 6038 2086
rect 6026 2076 6028 2084
rect 6036 2076 6038 2084
rect 6026 1824 6038 2076
rect 6090 2064 6102 2656
rect 6154 2704 6166 2706
rect 6154 2696 6156 2704
rect 6164 2696 6166 2704
rect 6090 2056 6092 2064
rect 6100 2056 6102 2064
rect 6090 2054 6102 2056
rect 6122 2644 6134 2646
rect 6122 2636 6124 2644
rect 6132 2636 6134 2644
rect 6026 1816 6028 1824
rect 6036 1816 6038 1824
rect 6026 1724 6038 1816
rect 6026 1716 6028 1724
rect 6036 1716 6038 1724
rect 6026 1424 6038 1716
rect 6090 2004 6102 2006
rect 6090 1996 6092 2004
rect 6100 1996 6102 2004
rect 6026 1416 6028 1424
rect 6036 1416 6038 1424
rect 6026 1414 6038 1416
rect 6058 1504 6070 1506
rect 6058 1496 6060 1504
rect 6068 1496 6070 1504
rect 5994 1336 5996 1344
rect 6004 1336 6006 1344
rect 5930 936 5932 944
rect 5940 936 5942 944
rect 5930 934 5942 936
rect 5962 1084 5974 1086
rect 5962 1076 5964 1084
rect 5972 1076 5974 1084
rect 5898 916 5900 924
rect 5908 916 5910 924
rect 5898 914 5910 916
rect 5930 904 5942 906
rect 5930 896 5932 904
rect 5940 896 5942 904
rect 5866 496 5868 504
rect 5876 496 5878 504
rect 5866 304 5878 496
rect 5866 296 5868 304
rect 5876 296 5878 304
rect 5866 294 5878 296
rect 5898 884 5910 886
rect 5898 876 5900 884
rect 5908 876 5910 884
rect 5898 184 5910 876
rect 5930 784 5942 896
rect 5962 844 5974 1076
rect 5994 1084 6006 1336
rect 5994 1076 5996 1084
rect 6004 1076 6006 1084
rect 5994 964 6006 1076
rect 5994 956 5996 964
rect 6004 956 6006 964
rect 5994 954 6006 956
rect 6026 1364 6038 1366
rect 6026 1356 6028 1364
rect 6036 1356 6038 1364
rect 5962 836 5964 844
rect 5972 836 5974 844
rect 5962 834 5974 836
rect 5994 864 6006 866
rect 5994 856 5996 864
rect 6004 856 6006 864
rect 5930 776 5932 784
rect 5940 776 5942 784
rect 5930 774 5942 776
rect 5962 784 5974 786
rect 5962 776 5964 784
rect 5972 776 5974 784
rect 5930 724 5942 726
rect 5930 716 5932 724
rect 5940 716 5942 724
rect 5930 404 5942 716
rect 5962 464 5974 776
rect 5994 684 6006 856
rect 5994 676 5996 684
rect 6004 676 6006 684
rect 5994 674 6006 676
rect 5962 456 5964 464
rect 5972 456 5974 464
rect 5962 454 5974 456
rect 5994 584 6006 586
rect 5994 576 5996 584
rect 6004 576 6006 584
rect 5930 396 5932 404
rect 5940 396 5942 404
rect 5930 394 5942 396
rect 5962 384 5974 386
rect 5962 376 5964 384
rect 5972 376 5974 384
rect 5930 364 5942 366
rect 5930 356 5932 364
rect 5940 356 5942 364
rect 5930 264 5942 356
rect 5962 304 5974 376
rect 5962 296 5964 304
rect 5972 296 5974 304
rect 5962 294 5974 296
rect 5930 256 5932 264
rect 5940 256 5942 264
rect 5930 254 5942 256
rect 5898 176 5900 184
rect 5908 176 5910 184
rect 5898 174 5910 176
rect 5930 184 5942 186
rect 5930 176 5932 184
rect 5940 176 5942 184
rect 5802 156 5804 164
rect 5812 156 5814 164
rect 5802 154 5814 156
rect 5738 116 5740 124
rect 5748 116 5750 124
rect 5738 114 5750 116
rect 5674 96 5676 104
rect 5684 96 5686 104
rect 5674 94 5686 96
rect 5930 84 5942 176
rect 5994 144 6006 576
rect 5994 136 5996 144
rect 6004 136 6006 144
rect 5994 134 6006 136
rect 6026 104 6038 1356
rect 6058 1284 6070 1496
rect 6058 1276 6060 1284
rect 6068 1276 6070 1284
rect 6058 1274 6070 1276
rect 6058 1224 6070 1226
rect 6058 1216 6060 1224
rect 6068 1216 6070 1224
rect 6058 784 6070 1216
rect 6058 776 6060 784
rect 6068 776 6070 784
rect 6058 774 6070 776
rect 6058 744 6070 746
rect 6058 736 6060 744
rect 6068 736 6070 744
rect 6058 324 6070 736
rect 6058 316 6060 324
rect 6068 316 6070 324
rect 6058 314 6070 316
rect 6090 524 6102 1996
rect 6122 944 6134 2636
rect 6154 2644 6166 2696
rect 6154 2636 6156 2644
rect 6164 2636 6166 2644
rect 6154 2634 6166 2636
rect 6186 2684 6198 2686
rect 6186 2676 6188 2684
rect 6196 2676 6198 2684
rect 6122 936 6124 944
rect 6132 936 6134 944
rect 6122 934 6134 936
rect 6154 2604 6166 2606
rect 6154 2596 6156 2604
rect 6164 2596 6166 2604
rect 6154 904 6166 2596
rect 6186 1124 6198 2676
rect 6218 1204 6230 4116
rect 6250 2544 6262 4336
rect 6282 4084 6294 4086
rect 6282 4076 6284 4084
rect 6292 4076 6294 4084
rect 6282 3764 6294 4076
rect 6282 3756 6284 3764
rect 6292 3756 6294 3764
rect 6282 3754 6294 3756
rect 6250 2536 6252 2544
rect 6260 2536 6262 2544
rect 6250 2534 6262 2536
rect 6282 3704 6294 3706
rect 6282 3696 6284 3704
rect 6292 3696 6294 3704
rect 6250 2364 6262 2366
rect 6250 2356 6252 2364
rect 6260 2356 6262 2364
rect 6250 1884 6262 2356
rect 6250 1876 6252 1884
rect 6260 1876 6262 1884
rect 6250 1874 6262 1876
rect 6250 1704 6262 1706
rect 6250 1696 6252 1704
rect 6260 1696 6262 1704
rect 6250 1544 6262 1696
rect 6250 1536 6252 1544
rect 6260 1536 6262 1544
rect 6250 1534 6262 1536
rect 6218 1196 6220 1204
rect 6228 1196 6230 1204
rect 6218 1194 6230 1196
rect 6250 1504 6262 1506
rect 6250 1496 6252 1504
rect 6260 1496 6262 1504
rect 6186 1116 6188 1124
rect 6196 1116 6198 1124
rect 6186 1114 6198 1116
rect 6218 1164 6230 1166
rect 6218 1156 6220 1164
rect 6228 1156 6230 1164
rect 6154 896 6156 904
rect 6164 896 6166 904
rect 6154 894 6166 896
rect 6186 1004 6198 1006
rect 6186 996 6188 1004
rect 6196 996 6198 1004
rect 6090 516 6092 524
rect 6100 516 6102 524
rect 6090 124 6102 516
rect 6090 116 6092 124
rect 6100 116 6102 124
rect 6090 114 6102 116
rect 6122 784 6134 786
rect 6122 776 6124 784
rect 6132 776 6134 784
rect 6026 96 6028 104
rect 6036 96 6038 104
rect 6026 94 6038 96
rect 5930 76 5932 84
rect 5940 76 5942 84
rect 5930 74 5942 76
rect 5482 16 5484 24
rect 5492 16 5494 24
rect 5482 14 5494 16
rect 5738 64 5750 66
rect 5738 56 5740 64
rect 5748 56 5750 64
rect 5738 24 5750 56
rect 5738 16 5740 24
rect 5748 16 5750 24
rect 5738 14 5750 16
rect 6122 24 6134 776
rect 6154 684 6166 686
rect 6154 676 6156 684
rect 6164 676 6166 684
rect 6154 364 6166 676
rect 6154 356 6156 364
rect 6164 356 6166 364
rect 6154 354 6166 356
rect 6154 204 6166 206
rect 6154 196 6156 204
rect 6164 196 6166 204
rect 6154 144 6166 196
rect 6154 136 6156 144
rect 6164 136 6166 144
rect 6154 134 6166 136
rect 6186 124 6198 996
rect 6218 684 6230 1156
rect 6250 988 6262 1496
rect 6250 980 6252 988
rect 6260 980 6262 988
rect 6250 974 6262 980
rect 6250 960 6262 966
rect 6250 952 6252 960
rect 6260 952 6262 960
rect 6250 864 6262 952
rect 6250 856 6252 864
rect 6260 856 6262 864
rect 6250 854 6262 856
rect 6218 676 6220 684
rect 6228 676 6230 684
rect 6218 674 6230 676
rect 6250 704 6262 706
rect 6250 696 6252 704
rect 6260 696 6262 704
rect 6250 644 6262 696
rect 6250 636 6252 644
rect 6260 636 6262 644
rect 6250 634 6262 636
rect 6282 604 6294 3696
rect 6282 596 6284 604
rect 6292 596 6294 604
rect 6282 594 6294 596
rect 6250 564 6262 566
rect 6250 556 6252 564
rect 6260 556 6262 564
rect 6250 164 6262 556
rect 6250 156 6252 164
rect 6260 156 6262 164
rect 6250 154 6262 156
rect 6186 116 6188 124
rect 6196 116 6198 124
rect 6186 114 6198 116
rect 6122 16 6124 24
rect 6132 16 6134 24
rect 6122 14 6134 16
rect 4664 6 4666 14
rect 4674 6 4678 14
rect 4686 6 4690 14
rect 4698 6 4702 14
rect 4710 6 4712 14
rect 4664 -40 4712 6
use NAND2X1  NAND2X1_28
timestamp 1522732896
transform -1 0 56 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1522732896
transform -1 0 120 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_20
timestamp 1522732896
transform -1 0 152 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_72
timestamp 1522732896
transform -1 0 344 0 -1 4610
box 0 0 192 200
use BUFX4  BUFX4_24
timestamp 1522732896
transform -1 0 408 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_69
timestamp 1522732896
transform 1 0 408 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_25
timestamp 1522732896
transform 1 0 600 0 -1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_31
timestamp 1522732896
transform -1 0 680 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_29
timestamp 1522732896
transform -1 0 744 0 -1 4610
box 0 0 64 200
use BUFX2  BUFX2_26
timestamp 1522732896
transform -1 0 792 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_74
timestamp 1522732896
transform 1 0 792 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_10
timestamp 1522732896
transform 1 0 984 0 -1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_14
timestamp 1522732896
transform 1 0 1016 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_8
timestamp 1522732896
transform 1 0 1064 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_12
timestamp 1522732896
transform -1 0 1160 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_98
timestamp 1522732896
transform -1 0 1352 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_19
timestamp 1522732896
transform -1 0 1384 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_96
timestamp 1522732896
transform -1 0 1576 0 -1 4610
box 0 0 192 200
use FILL  FILL_22_0_0
timestamp 1522732896
transform 1 0 1576 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_1
timestamp 1522732896
transform 1 0 1592 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_2
timestamp 1522732896
transform 1 0 1608 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_324
timestamp 1522732896
transform 1 0 1624 0 -1 4610
box 0 0 64 200
use BUFX2  BUFX2_22
timestamp 1522732896
transform 1 0 1688 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_323
timestamp 1522732896
transform -1 0 1800 0 -1 4610
box 0 0 64 200
use OR2X2  OR2X2_30
timestamp 1522732896
transform 1 0 1800 0 -1 4610
box 0 0 64 200
use BUFX2  BUFX2_19
timestamp 1522732896
transform 1 0 1864 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_23
timestamp 1522732896
transform 1 0 1912 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_30
timestamp 1522732896
transform -1 0 2008 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_32
timestamp 1522732896
transform -1 0 2056 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_20
timestamp 1522732896
transform 1 0 2056 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1522732896
transform 1 0 2104 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_237
timestamp 1522732896
transform 1 0 2296 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_169
timestamp 1522732896
transform -1 0 2408 0 -1 4610
box 0 0 48 200
use INVX1  INVX1_82
timestamp 1522732896
transform -1 0 2440 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1522732896
transform -1 0 2632 0 -1 4610
box 0 0 192 200
use BUFX2  BUFX2_35
timestamp 1522732896
transform -1 0 2680 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_183
timestamp 1522732896
transform 1 0 2680 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_285
timestamp 1522732896
transform -1 0 2792 0 -1 4610
box 0 0 64 200
use BUFX2  BUFX2_40
timestamp 1522732896
transform -1 0 2840 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1522732896
transform 1 0 2840 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_100
timestamp 1522732896
transform 1 0 3032 0 -1 4610
box 0 0 32 200
use BUFX2  BUFX2_36
timestamp 1522732896
transform -1 0 3112 0 -1 4610
box 0 0 48 200
use FILL  FILL_22_1_0
timestamp 1522732896
transform -1 0 3128 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_1
timestamp 1522732896
transform -1 0 3144 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_2
timestamp 1522732896
transform -1 0 3160 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1522732896
transform -1 0 3352 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_290
timestamp 1522732896
transform 1 0 3352 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_188
timestamp 1522732896
transform -1 0 3464 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1522732896
transform 1 0 3464 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_92
timestamp 1522732896
transform -1 0 3688 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1522732896
transform -1 0 3880 0 -1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1522732896
transform 1 0 3880 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_99
timestamp 1522732896
transform -1 0 4104 0 -1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_187
timestamp 1522732896
transform 1 0 4104 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_289
timestamp 1522732896
transform -1 0 4216 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1522732896
transform -1 0 4408 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_96
timestamp 1522732896
transform -1 0 4440 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1522732896
transform -1 0 4632 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_97
timestamp 1522732896
transform -1 0 4664 0 -1 4610
box 0 0 32 200
use FILL  FILL_22_2_0
timestamp 1522732896
transform 1 0 4664 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_1
timestamp 1522732896
transform 1 0 4680 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_2
timestamp 1522732896
transform 1 0 4696 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_241
timestamp 1522732896
transform 1 0 4712 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_173
timestamp 1522732896
transform -1 0 4824 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1522732896
transform -1 0 5016 0 -1 4610
box 0 0 192 200
use BUFX4  BUFX4_18
timestamp 1522732896
transform 1 0 5016 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_244
timestamp 1522732896
transform 1 0 5080 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_129
timestamp 1522732896
transform -1 0 5320 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_463
timestamp 1522732896
transform -1 0 5384 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_433
timestamp 1522732896
transform -1 0 5448 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_229
timestamp 1522732896
transform -1 0 5496 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_228
timestamp 1522732896
transform -1 0 5544 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_235
timestamp 1522732896
transform 1 0 5544 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_172
timestamp 1522732896
transform 1 0 5592 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_168
timestamp 1522732896
transform -1 0 5720 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_171
timestamp 1522732896
transform 1 0 5720 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_227
timestamp 1522732896
transform -1 0 5832 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_226
timestamp 1522732896
transform -1 0 5880 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_462
timestamp 1522732896
transform -1 0 5944 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_225
timestamp 1522732896
transform 1 0 5944 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_429
timestamp 1522732896
transform 1 0 5992 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_236
timestamp 1522732896
transform -1 0 6104 0 -1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_37
timestamp 1522732896
transform -1 0 6184 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_461
timestamp 1522732896
transform 1 0 6184 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_252
timestamp 1522732896
transform -1 0 6296 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_121
timestamp 1522732896
transform -1 0 200 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_94
timestamp 1522732896
transform 1 0 200 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_101
timestamp 1522732896
transform 1 0 392 0 1 4210
box 0 0 192 200
use BUFX2  BUFX2_17
timestamp 1522732896
transform -1 0 632 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_104
timestamp 1522732896
transform 1 0 632 0 1 4210
box 0 0 192 200
use OR2X2  OR2X2_26
timestamp 1522732896
transform -1 0 888 0 1 4210
box 0 0 64 200
use BUFX2  BUFX2_24
timestamp 1522732896
transform -1 0 936 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_332
timestamp 1522732896
transform -1 0 1000 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_331
timestamp 1522732896
transform -1 0 1064 0 1 4210
box 0 0 64 200
use OR2X2  OR2X2_32
timestamp 1522732896
transform 1 0 1064 0 1 4210
box 0 0 64 200
use BUFX2  BUFX2_21
timestamp 1522732896
transform 1 0 1128 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_97
timestamp 1522732896
transform 1 0 1176 0 1 4210
box 0 0 192 200
use BUFX2  BUFX2_27
timestamp 1522732896
transform 1 0 1368 0 1 4210
box 0 0 48 200
use OR2X2  OR2X2_34
timestamp 1522732896
transform -1 0 1480 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_339
timestamp 1522732896
transform 1 0 1480 0 1 4210
box 0 0 64 200
use BUFX2  BUFX2_31
timestamp 1522732896
transform 1 0 1544 0 1 4210
box 0 0 48 200
use FILL  FILL_21_0_0
timestamp 1522732896
transform 1 0 1592 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_1
timestamp 1522732896
transform 1 0 1608 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_2
timestamp 1522732896
transform 1 0 1624 0 1 4210
box 0 0 16 200
use BUFX2  BUFX2_29
timestamp 1522732896
transform 1 0 1640 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1522732896
transform -1 0 1880 0 1 4210
box 0 0 192 200
use INVX1  INVX1_81
timestamp 1522732896
transform 1 0 1880 0 1 4210
box 0 0 32 200
use MUX2X1  MUX2X1_29
timestamp 1522732896
transform -1 0 2008 0 1 4210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1522732896
transform 1 0 2008 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_174
timestamp 1522732896
transform 1 0 2200 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_242
timestamp 1522732896
transform -1 0 2312 0 1 4210
box 0 0 64 200
use INVX1  INVX1_101
timestamp 1522732896
transform 1 0 2312 0 1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_140
timestamp 1522732896
transform 1 0 2344 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_131
timestamp 1522732896
transform 1 0 2392 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1522732896
transform 1 0 2440 0 1 4210
box 0 0 192 200
use INVX1  INVX1_79
timestamp 1522732896
transform 1 0 2632 0 1 4210
box 0 0 32 200
use MUX2X1  MUX2X1_13
timestamp 1522732896
transform -1 0 2760 0 1 4210
box 0 0 96 200
use MUX2X1  MUX2X1_20
timestamp 1522732896
transform -1 0 2856 0 1 4210
box 0 0 96 200
use BUFX2  BUFX2_39
timestamp 1522732896
transform 1 0 2856 0 1 4210
box 0 0 48 200
use MUX2X1  MUX2X1_34
timestamp 1522732896
transform -1 0 3000 0 1 4210
box 0 0 96 200
use INVX1  INVX1_102
timestamp 1522732896
transform -1 0 3032 0 1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_141
timestamp 1522732896
transform -1 0 3080 0 1 4210
box 0 0 48 200
use INVX1  INVX1_103
timestamp 1522732896
transform -1 0 3112 0 1 4210
box 0 0 32 200
use FILL  FILL_21_1_0
timestamp 1522732896
transform 1 0 3112 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_1
timestamp 1522732896
transform 1 0 3128 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_2
timestamp 1522732896
transform 1 0 3144 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1522732896
transform 1 0 3160 0 1 4210
box 0 0 192 200
use INVX1  INVX1_94
timestamp 1522732896
transform 1 0 3352 0 1 4210
box 0 0 32 200
use MUX2X1  MUX2X1_32
timestamp 1522732896
transform 1 0 3384 0 1 4210
box 0 0 96 200
use MUX2X1  MUX2X1_17
timestamp 1522732896
transform -1 0 3576 0 1 4210
box 0 0 96 200
use OAI21X1  OAI21X1_240
timestamp 1522732896
transform 1 0 3576 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_172
timestamp 1522732896
transform -1 0 3688 0 1 4210
box 0 0 48 200
use INVX1  INVX1_93
timestamp 1522732896
transform 1 0 3688 0 1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_136
timestamp 1522732896
transform 1 0 3720 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1522732896
transform -1 0 3960 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_139
timestamp 1522732896
transform -1 0 4008 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1522732896
transform 1 0 4008 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_138
timestamp 1522732896
transform -1 0 4248 0 1 4210
box 0 0 48 200
use INVX1  INVX1_98
timestamp 1522732896
transform 1 0 4248 0 1 4210
box 0 0 32 200
use MUX2X1  MUX2X1_33
timestamp 1522732896
transform 1 0 4280 0 1 4210
box 0 0 96 200
use MUX2X1  MUX2X1_18
timestamp 1522732896
transform 1 0 4376 0 1 4210
box 0 0 96 200
use NAND2X1  NAND2X1_167
timestamp 1522732896
transform 1 0 4472 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_235
timestamp 1522732896
transform -1 0 4584 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_283
timestamp 1522732896
transform 1 0 4584 0 1 4210
box 0 0 64 200
use FILL  FILL_21_2_0
timestamp 1522732896
transform -1 0 4664 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_1
timestamp 1522732896
transform -1 0 4680 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_2
timestamp 1522732896
transform -1 0 4696 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_181
timestamp 1522732896
transform -1 0 4744 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1522732896
transform -1 0 4936 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_131
timestamp 1522732896
transform -1 0 5128 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_246
timestamp 1522732896
transform 1 0 5128 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_465
timestamp 1522732896
transform -1 0 5240 0 1 4210
box 0 0 64 200
use XNOR2X1  XNOR2X1_8
timestamp 1522732896
transform -1 0 5352 0 1 4210
box 0 0 112 200
use OAI21X1  OAI21X1_432
timestamp 1522732896
transform 1 0 5352 0 1 4210
box 0 0 64 200
use INVX1  INVX1_184
timestamp 1522732896
transform -1 0 5448 0 1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_124
timestamp 1522732896
transform 1 0 5448 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_56
timestamp 1522732896
transform -1 0 5592 0 1 4210
box 0 0 80 200
use MUX2X1  MUX2X1_36
timestamp 1522732896
transform 1 0 5592 0 1 4210
box 0 0 96 200
use OAI21X1  OAI21X1_410
timestamp 1522732896
transform -1 0 5752 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_421
timestamp 1522732896
transform -1 0 5816 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_431
timestamp 1522732896
transform -1 0 5880 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_414
timestamp 1522732896
transform -1 0 5944 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_234
timestamp 1522732896
transform -1 0 5992 0 1 4210
box 0 0 48 200
use INVX1  INVX1_177
timestamp 1522732896
transform -1 0 6024 0 1 4210
box 0 0 32 200
use INVX1  INVX1_183
timestamp 1522732896
transform -1 0 6056 0 1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_131
timestamp 1522732896
transform -1 0 6120 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_428
timestamp 1522732896
transform -1 0 6184 0 1 4210
box 0 0 64 200
use INVX1  INVX1_182
timestamp 1522732896
transform 1 0 6184 0 1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_228
timestamp 1522732896
transform -1 0 6264 0 1 4210
box 0 0 48 200
use FILL  FILL_22_1
timestamp 1522732896
transform 1 0 6264 0 1 4210
box 0 0 16 200
use FILL  FILL_22_2
timestamp 1522732896
transform 1 0 6280 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_120
timestamp 1522732896
transform 1 0 8 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_391
timestamp 1522732896
transform -1 0 264 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_161
timestamp 1522732896
transform -1 0 296 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_222
timestamp 1522732896
transform -1 0 344 0 -1 4210
box 0 0 48 200
use OAI22X1  OAI22X1_52
timestamp 1522732896
transform -1 0 424 0 -1 4210
box 0 0 80 200
use INVX2  INVX2_17
timestamp 1522732896
transform 1 0 424 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_114
timestamp 1522732896
transform 1 0 456 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_13
timestamp 1522732896
transform 1 0 648 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_99
timestamp 1522732896
transform 1 0 680 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_11
timestamp 1522732896
transform 1 0 872 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_344
timestamp 1522732896
transform 1 0 904 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_336
timestamp 1522732896
transform 1 0 968 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_315
timestamp 1522732896
transform 1 0 1032 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_316
timestamp 1522732896
transform -1 0 1160 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_152
timestamp 1522732896
transform -1 0 1192 0 -1 4210
box 0 0 32 200
use BUFX4  BUFX4_55
timestamp 1522732896
transform -1 0 1256 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_356
timestamp 1522732896
transform -1 0 1320 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_17
timestamp 1522732896
transform 1 0 1320 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_199
timestamp 1522732896
transform -1 0 1400 0 -1 4210
box 0 0 48 200
use OR2X2  OR2X2_35
timestamp 1522732896
transform -1 0 1464 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_343
timestamp 1522732896
transform -1 0 1528 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_56
timestamp 1522732896
transform -1 0 1592 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_0_0
timestamp 1522732896
transform -1 0 1608 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_1
timestamp 1522732896
transform -1 0 1624 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_2
timestamp 1522732896
transform -1 0 1640 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_335
timestamp 1522732896
transform -1 0 1704 0 -1 4210
box 0 0 64 200
use OR2X2  OR2X2_33
timestamp 1522732896
transform -1 0 1768 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_328
timestamp 1522732896
transform 1 0 1768 0 -1 4210
box 0 0 64 200
use BUFX2  BUFX2_18
timestamp 1522732896
transform -1 0 1880 0 -1 4210
box 0 0 48 200
use BUFX4  BUFX4_57
timestamp 1522732896
transform 1 0 1880 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_340
timestamp 1522732896
transform -1 0 2008 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_14
timestamp 1522732896
transform -1 0 2040 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_100
timestamp 1522732896
transform -1 0 2232 0 -1 4210
box 0 0 192 200
use BUFX4  BUFX4_15
timestamp 1522732896
transform -1 0 2296 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_34
timestamp 1522732896
transform -1 0 2488 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_80
timestamp 1522732896
transform 1 0 2488 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_130
timestamp 1522732896
transform 1 0 2520 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_110
timestamp 1522732896
transform -1 0 2632 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_108
timestamp 1522732896
transform -1 0 2696 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_109
timestamp 1522732896
transform 1 0 2696 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_107
timestamp 1522732896
transform 1 0 2760 0 -1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_105
timestamp 1522732896
transform -1 0 2888 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_128
timestamp 1522732896
transform 1 0 2888 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_127
timestamp 1522732896
transform 1 0 2952 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_130
timestamp 1522732896
transform 1 0 3016 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_129
timestamp 1522732896
transform 1 0 3080 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_1_0
timestamp 1522732896
transform -1 0 3160 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_1
timestamp 1522732896
transform -1 0 3176 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_2
timestamp 1522732896
transform -1 0 3192 0 -1 4210
box 0 0 16 200
use AOI21X1  AOI21X1_103
timestamp 1522732896
transform -1 0 3256 0 -1 4210
box 0 0 64 200
use BUFX2  BUFX2_38
timestamp 1522732896
transform 1 0 3256 0 -1 4210
box 0 0 48 200
use AOI21X1  AOI21X1_101
timestamp 1522732896
transform -1 0 3368 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1522732896
transform 1 0 3368 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_85
timestamp 1522732896
transform 1 0 3560 0 -1 4210
box 0 0 32 200
use MUX2X1  MUX2X1_30
timestamp 1522732896
transform 1 0 3592 0 -1 4210
box 0 0 96 200
use NAND3X1  NAND3X1_113
timestamp 1522732896
transform 1 0 3688 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_120
timestamp 1522732896
transform 1 0 3752 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_119
timestamp 1522732896
transform 1 0 3816 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_111
timestamp 1522732896
transform -1 0 3944 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_126
timestamp 1522732896
transform 1 0 3944 0 -1 4210
box 0 0 64 200
use MUX2X1  MUX2X1_15
timestamp 1522732896
transform 1 0 4008 0 -1 4210
box 0 0 96 200
use INVX1  INVX1_83
timestamp 1522732896
transform -1 0 4136 0 -1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_124
timestamp 1522732896
transform 1 0 4136 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_125
timestamp 1522732896
transform -1 0 4264 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_99
timestamp 1522732896
transform -1 0 4328 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_123
timestamp 1522732896
transform -1 0 4392 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_71
timestamp 1522732896
transform -1 0 4424 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1522732896
transform -1 0 4616 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_73
timestamp 1522732896
transform -1 0 4648 0 -1 4210
box 0 0 32 200
use FILL  FILL_20_2_0
timestamp 1522732896
transform 1 0 4648 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_1
timestamp 1522732896
transform 1 0 4664 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_2
timestamp 1522732896
transform 1 0 4680 0 -1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_27
timestamp 1522732896
transform 1 0 4696 0 -1 4210
box 0 0 96 200
use INVX1  INVX1_72
timestamp 1522732896
transform -1 0 4824 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1522732896
transform -1 0 5016 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_466
timestamp 1522732896
transform -1 0 5080 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_181
timestamp 1522732896
transform 1 0 5080 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_236
timestamp 1522732896
transform 1 0 5112 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_456
timestamp 1522732896
transform 1 0 5160 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_427
timestamp 1522732896
transform 1 0 5224 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_426
timestamp 1522732896
transform -1 0 5352 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_434
timestamp 1522732896
transform -1 0 5416 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_201
timestamp 1522732896
transform -1 0 5448 0 -1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_125
timestamp 1522732896
transform -1 0 5512 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_232
timestamp 1522732896
transform -1 0 5560 0 -1 4210
box 0 0 48 200
use XOR2X1  XOR2X1_2
timestamp 1522732896
transform -1 0 5672 0 -1 4210
box 0 0 112 200
use OAI21X1  OAI21X1_409
timestamp 1522732896
transform 1 0 5672 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_408
timestamp 1522732896
transform -1 0 5800 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_412
timestamp 1522732896
transform 1 0 5800 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_413
timestamp 1522732896
transform -1 0 5928 0 -1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_123
timestamp 1522732896
transform -1 0 5992 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_430
timestamp 1522732896
transform -1 0 6056 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_55
timestamp 1522732896
transform -1 0 6136 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_418
timestamp 1522732896
transform -1 0 6200 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_167
timestamp 1522732896
transform 1 0 6200 0 -1 4210
box 0 0 64 200
use FILL  FILL_21_1
timestamp 1522732896
transform -1 0 6280 0 -1 4210
box 0 0 16 200
use FILL  FILL_21_2
timestamp 1522732896
transform -1 0 6296 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_160
timestamp 1522732896
transform 1 0 8 0 1 3810
box 0 0 32 200
use NOR2X1  NOR2X1_221
timestamp 1522732896
transform 1 0 40 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_393
timestamp 1522732896
transform -1 0 152 0 1 3810
box 0 0 64 200
use OAI22X1  OAI22X1_53
timestamp 1522732896
transform -1 0 232 0 1 3810
box 0 0 80 200
use INVX2  INVX2_15
timestamp 1522732896
transform 1 0 232 0 1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_120
timestamp 1522732896
transform 1 0 264 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_392
timestamp 1522732896
transform 1 0 328 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_390
timestamp 1522732896
transform 1 0 392 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_380
timestamp 1522732896
transform -1 0 520 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_26
timestamp 1522732896
transform 1 0 520 0 1 3810
box 0 0 64 200
use INVX2  INVX2_5
timestamp 1522732896
transform -1 0 616 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_103
timestamp 1522732896
transform 1 0 616 0 1 3810
box 0 0 192 200
use INVX1  INVX1_24
timestamp 1522732896
transform 1 0 808 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_352
timestamp 1522732896
transform 1 0 840 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_198
timestamp 1522732896
transform -1 0 952 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_17
timestamp 1522732896
transform -1 0 1016 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1522732896
transform 1 0 1016 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_312
timestamp 1522732896
transform 1 0 1080 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_15
timestamp 1522732896
transform 1 0 1144 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_311
timestamp 1522732896
transform 1 0 1208 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_90
timestamp 1522732896
transform -1 0 1336 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_330
timestamp 1522732896
transform 1 0 1336 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_333
timestamp 1522732896
transform 1 0 1400 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_102
timestamp 1522732896
transform -1 0 1528 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_334
timestamp 1522732896
transform -1 0 1592 0 1 3810
box 0 0 64 200
use FILL  FILL_19_0_0
timestamp 1522732896
transform 1 0 1592 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1522732896
transform 1 0 1608 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_2
timestamp 1522732896
transform 1 0 1624 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_321
timestamp 1522732896
transform 1 0 1640 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_96
timestamp 1522732896
transform -1 0 1768 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_322
timestamp 1522732896
transform -1 0 1832 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_325
timestamp 1522732896
transform 1 0 1832 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_98
timestamp 1522732896
transform -1 0 1960 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_327
timestamp 1522732896
transform -1 0 2024 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_326
timestamp 1522732896
transform -1 0 2088 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_31
timestamp 1522732896
transform 1 0 2088 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_28
timestamp 1522732896
transform -1 0 2200 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_25
timestamp 1522732896
transform 1 0 2200 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_89
timestamp 1522732896
transform -1 0 2312 0 1 3810
box 0 0 64 200
use INVX1  INVX1_129
timestamp 1522732896
transform 1 0 2312 0 1 3810
box 0 0 32 200
use NAND3X1  NAND3X1_135
timestamp 1522732896
transform -1 0 2408 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_26
timestamp 1522732896
transform 1 0 2408 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_33
timestamp 1522732896
transform 1 0 2472 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_95
timestamp 1522732896
transform -1 0 2584 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_29
timestamp 1522732896
transform 1 0 2584 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_43
timestamp 1522732896
transform 1 0 2648 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_166
timestamp 1522732896
transform 1 0 2712 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_131
timestamp 1522732896
transform -1 0 2824 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_192
timestamp 1522732896
transform 1 0 2824 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_153
timestamp 1522732896
transform -1 0 2920 0 1 3810
box 0 0 48 200
use AND2X2  AND2X2_34
timestamp 1522732896
transform 1 0 2920 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_47
timestamp 1522732896
transform -1 0 3048 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_97
timestamp 1522732896
transform -1 0 3112 0 1 3810
box 0 0 64 200
use FILL  FILL_19_1_0
timestamp 1522732896
transform 1 0 3112 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1522732896
transform 1 0 3128 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_2
timestamp 1522732896
transform 1 0 3144 0 1 3810
box 0 0 16 200
use AND2X2  AND2X2_30
timestamp 1522732896
transform 1 0 3160 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_33
timestamp 1522732896
transform -1 0 3288 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_2
timestamp 1522732896
transform -1 0 3336 0 1 3810
box 0 0 48 200
use AND2X2  AND2X2_32
timestamp 1522732896
transform -1 0 3400 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_77
timestamp 1522732896
transform -1 0 3464 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_122
timestamp 1522732896
transform 1 0 3464 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_121
timestamp 1522732896
transform 1 0 3528 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_6
timestamp 1522732896
transform -1 0 3640 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_14
timestamp 1522732896
transform -1 0 3688 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_114
timestamp 1522732896
transform -1 0 3752 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_112
timestamp 1522732896
transform 1 0 3752 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_137
timestamp 1522732896
transform -1 0 3864 0 1 3810
box 0 0 48 200
use INVX1  INVX1_95
timestamp 1522732896
transform -1 0 3896 0 1 3810
box 0 0 32 200
use BUFX2  BUFX2_3
timestamp 1522732896
transform -1 0 3944 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_98
timestamp 1522732896
transform 1 0 3944 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_126
timestamp 1522732896
transform -1 0 4056 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_100
timestamp 1522732896
transform 1 0 4056 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_127
timestamp 1522732896
transform -1 0 4168 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_13
timestamp 1522732896
transform 1 0 4168 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_97
timestamp 1522732896
transform -1 0 4280 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_288
timestamp 1522732896
transform 1 0 4280 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_186
timestamp 1522732896
transform -1 0 4392 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1522732896
transform -1 0 4584 0 1 3810
box 0 0 192 200
use FILL  FILL_19_2_0
timestamp 1522732896
transform -1 0 4600 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1522732896
transform -1 0 4616 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_2
timestamp 1522732896
transform -1 0 4632 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_133
timestamp 1522732896
transform -1 0 4824 0 1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_132
timestamp 1522732896
transform -1 0 5016 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_247
timestamp 1522732896
transform 1 0 5016 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_468
timestamp 1522732896
transform -1 0 5128 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_467
timestamp 1522732896
transform -1 0 5192 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_239
timestamp 1522732896
transform -1 0 5240 0 1 3810
box 0 0 48 200
use INVX1  INVX1_204
timestamp 1522732896
transform 1 0 5240 0 1 3810
box 0 0 32 200
use AOI22X1  AOI22X1_62
timestamp 1522732896
transform -1 0 5352 0 1 3810
box 0 0 80 200
use INVX1  INVX1_168
timestamp 1522732896
transform -1 0 5384 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_455
timestamp 1522732896
transform 1 0 5384 0 1 3810
box 0 0 64 200
use INVX1  INVX1_202
timestamp 1522732896
transform 1 0 5448 0 1 3810
box 0 0 32 200
use AOI22X1  AOI22X1_60
timestamp 1522732896
transform -1 0 5560 0 1 3810
box 0 0 80 200
use OR2X2  OR2X2_40
timestamp 1522732896
transform -1 0 5624 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_233
timestamp 1522732896
transform -1 0 5672 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_451
timestamp 1522732896
transform -1 0 5736 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_420
timestamp 1522732896
transform -1 0 5800 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_231
timestamp 1522732896
transform -1 0 5848 0 1 3810
box 0 0 48 200
use INVX2  INVX2_45
timestamp 1522732896
transform -1 0 5880 0 1 3810
box 0 0 32 200
use NOR2X1  NOR2X1_233
timestamp 1522732896
transform -1 0 5928 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_417
timestamp 1522732896
transform 1 0 5928 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_416
timestamp 1522732896
transform -1 0 6056 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_54
timestamp 1522732896
transform -1 0 6136 0 1 3810
box 0 0 80 200
use AOI21X1  AOI21X1_122
timestamp 1522732896
transform -1 0 6200 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_222
timestamp 1522732896
transform 1 0 6200 0 1 3810
box 0 0 48 200
use FILL  FILL_20_1
timestamp 1522732896
transform 1 0 6248 0 1 3810
box 0 0 16 200
use FILL  FILL_20_2
timestamp 1522732896
transform 1 0 6264 0 1 3810
box 0 0 16 200
use FILL  FILL_20_3
timestamp 1522732896
transform 1 0 6280 0 1 3810
box 0 0 16 200
use OR2X2  OR2X2_37
timestamp 1522732896
transform -1 0 72 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_389
timestamp 1522732896
transform 1 0 72 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_211
timestamp 1522732896
transform 1 0 136 0 -1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_119
timestamp 1522732896
transform 1 0 184 0 -1 3810
box 0 0 64 200
use OAI22X1  OAI22X1_51
timestamp 1522732896
transform -1 0 328 0 -1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_33
timestamp 1522732896
transform -1 0 376 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_29
timestamp 1522732896
transform -1 0 440 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_9
timestamp 1522732896
transform -1 0 520 0 -1 3810
box 0 0 80 200
use NAND3X1  NAND3X1_26
timestamp 1522732896
transform 1 0 520 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_388
timestamp 1522732896
transform 1 0 584 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_119
timestamp 1522732896
transform 1 0 648 0 -1 3810
box 0 0 192 200
use INVX2  INVX2_18
timestamp 1522732896
transform -1 0 872 0 -1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_21
timestamp 1522732896
transform 1 0 872 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_23
timestamp 1522732896
transform -1 0 1000 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_29
timestamp 1522732896
transform -1 0 1048 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_28
timestamp 1522732896
transform 1 0 1048 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_32
timestamp 1522732896
transform 1 0 1112 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_22
timestamp 1522732896
transform -1 0 1224 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_27
timestamp 1522732896
transform -1 0 1272 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_351
timestamp 1522732896
transform 1 0 1272 0 -1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_6
timestamp 1522732896
transform -1 0 1400 0 -1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_24
timestamp 1522732896
transform 1 0 1400 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_43
timestamp 1522732896
transform -1 0 1544 0 -1 3810
box 0 0 80 200
use AOI22X1  AOI22X1_48
timestamp 1522732896
transform -1 0 1624 0 -1 3810
box 0 0 80 200
use FILL  FILL_18_0_0
timestamp 1522732896
transform 1 0 1624 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1522732896
transform 1 0 1640 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_2
timestamp 1522732896
transform 1 0 1656 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_329
timestamp 1522732896
transform 1 0 1672 0 -1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_100
timestamp 1522732896
transform -1 0 1800 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_45
timestamp 1522732896
transform -1 0 1880 0 -1 3810
box 0 0 80 200
use AOI22X1  AOI22X1_46
timestamp 1522732896
transform -1 0 1960 0 -1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_355
timestamp 1522732896
transform 1 0 1960 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1522732896
transform 1 0 2024 0 -1 3810
box 0 0 32 200
use BUFX4  BUFX4_53
timestamp 1522732896
transform 1 0 2056 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_200
timestamp 1522732896
transform -1 0 2168 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_105
timestamp 1522732896
transform 1 0 2168 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_359
timestamp 1522732896
transform 1 0 2360 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_167
timestamp 1522732896
transform -1 0 2488 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_71
timestamp 1522732896
transform 1 0 2488 0 -1 3810
box 0 0 192 200
use MUX2X1  MUX2X1_1
timestamp 1522732896
transform 1 0 2680 0 -1 3810
box 0 0 96 200
use NAND2X1  NAND2X1_180
timestamp 1522732896
transform -1 0 2824 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_172
timestamp 1522732896
transform -1 0 2888 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_155
timestamp 1522732896
transform -1 0 2952 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_182
timestamp 1522732896
transform 1 0 2952 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_180
timestamp 1522732896
transform -1 0 3080 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_174
timestamp 1522732896
transform -1 0 3144 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_1_0
timestamp 1522732896
transform -1 0 3160 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1522732896
transform -1 0 3176 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_2
timestamp 1522732896
transform -1 0 3192 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_156
timestamp 1522732896
transform -1 0 3256 0 -1 3810
box 0 0 64 200
use BUFX2  BUFX2_37
timestamp 1522732896
transform -1 0 3304 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_178
timestamp 1522732896
transform -1 0 3368 0 -1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_99
timestamp 1522732896
transform -1 0 3432 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1522732896
transform 1 0 3432 0 -1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_170
timestamp 1522732896
transform 1 0 3624 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_238
timestamp 1522732896
transform -1 0 3736 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_84
timestamp 1522732896
transform 1 0 3736 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_132
timestamp 1522732896
transform 1 0 3768 0 -1 3810
box 0 0 48 200
use BUFX4  BUFX4_46
timestamp 1522732896
transform 1 0 3816 0 -1 3810
box 0 0 64 200
use BUFX2  BUFX2_1
timestamp 1522732896
transform -1 0 3928 0 -1 3810
box 0 0 48 200
use BUFX2  BUFX2_15
timestamp 1522732896
transform 1 0 3928 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_106
timestamp 1522732896
transform 1 0 3976 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_105
timestamp 1522732896
transform -1 0 4104 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_117
timestamp 1522732896
transform -1 0 4168 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_129
timestamp 1522732896
transform -1 0 4216 0 -1 3810
box 0 0 48 200
use MUX2X1  MUX2X1_31
timestamp 1522732896
transform 1 0 4216 0 -1 3810
box 0 0 96 200
use INVX1  INVX1_89
timestamp 1522732896
transform -1 0 4344 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1522732896
transform -1 0 4536 0 -1 3810
box 0 0 192 200
use MUX2X1  MUX2X1_28
timestamp 1522732896
transform 1 0 4536 0 -1 3810
box 0 0 96 200
use INVX1  INVX1_77
timestamp 1522732896
transform -1 0 4664 0 -1 3810
box 0 0 32 200
use FILL  FILL_18_2_0
timestamp 1522732896
transform -1 0 4680 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1522732896
transform -1 0 4696 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_2
timestamp 1522732896
transform -1 0 4712 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1522732896
transform -1 0 4904 0 -1 3810
box 0 0 192 200
use BUFX4  BUFX4_21
timestamp 1522732896
transform 1 0 4904 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_248
timestamp 1522732896
transform 1 0 4968 0 -1 3810
box 0 0 48 200
use INVX8  INVX8_7
timestamp 1522732896
transform -1 0 5096 0 -1 3810
box 0 0 80 200
use BUFX4  BUFX4_65
timestamp 1522732896
transform -1 0 5160 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_172
timestamp 1522732896
transform 1 0 5160 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_425
timestamp 1522732896
transform -1 0 5256 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_49
timestamp 1522732896
transform -1 0 5320 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_424
timestamp 1522732896
transform -1 0 5384 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_407
timestamp 1522732896
transform 1 0 5384 0 -1 3810
box 0 0 64 200
use INVX2  INVX2_46
timestamp 1522732896
transform -1 0 5480 0 -1 3810
box 0 0 32 200
use INVX1  INVX1_174
timestamp 1522732896
transform 1 0 5480 0 -1 3810
box 0 0 32 200
use NAND3X1  NAND3X1_165
timestamp 1522732896
transform 1 0 5512 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_406
timestamp 1522732896
transform -1 0 5640 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_173
timestamp 1522732896
transform -1 0 5672 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_213
timestamp 1522732896
transform -1 0 5720 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_203
timestamp 1522732896
transform 1 0 5720 0 -1 3810
box 0 0 32 200
use AOI22X1  AOI22X1_53
timestamp 1522732896
transform 1 0 5752 0 -1 3810
box 0 0 80 200
use OAI22X1  OAI22X1_56
timestamp 1522732896
transform 1 0 5832 0 -1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_215
timestamp 1522732896
transform 1 0 5912 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_216
timestamp 1522732896
transform 1 0 5960 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_219
timestamp 1522732896
transform 1 0 6008 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_217
timestamp 1522732896
transform 1 0 6056 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_415
timestamp 1522732896
transform 1 0 6104 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_179
timestamp 1522732896
transform -1 0 6200 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_220
timestamp 1522732896
transform 1 0 6200 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_221
timestamp 1522732896
transform -1 0 6296 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_163
timestamp 1522732896
transform -1 0 72 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_387
timestamp 1522732896
transform -1 0 136 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_220
timestamp 1522732896
transform 1 0 136 0 1 3410
box 0 0 48 200
use AND2X2  AND2X2_47
timestamp 1522732896
transform 1 0 184 0 1 3410
box 0 0 64 200
use NOR3X1  NOR3X1_4
timestamp 1522732896
transform -1 0 376 0 1 3410
box 0 0 128 200
use INVX2  INVX2_19
timestamp 1522732896
transform -1 0 408 0 1 3410
box 0 0 32 200
use AND2X2  AND2X2_7
timestamp 1522732896
transform 1 0 408 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_386
timestamp 1522732896
transform 1 0 472 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_34
timestamp 1522732896
transform -1 0 600 0 1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_10
timestamp 1522732896
transform -1 0 680 0 1 3410
box 0 0 80 200
use AOI21X1  AOI21X1_27
timestamp 1522732896
transform 1 0 680 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1522732896
transform -1 0 808 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_30
timestamp 1522732896
transform 1 0 808 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_33
timestamp 1522732896
transform -1 0 936 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_19
timestamp 1522732896
transform 1 0 936 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_11
timestamp 1522732896
transform -1 0 1048 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1522732896
transform 1 0 1048 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_30
timestamp 1522732896
transform -1 0 1160 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_28
timestamp 1522732896
transform 1 0 1160 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1522732896
transform 1 0 1224 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_23
timestamp 1522732896
transform 1 0 1288 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1522732896
transform 1 0 1352 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_31
timestamp 1522732896
transform 1 0 1416 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_30
timestamp 1522732896
transform 1 0 1464 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_22
timestamp 1522732896
transform -1 0 1592 0 1 3410
box 0 0 64 200
use FILL  FILL_17_0_0
timestamp 1522732896
transform 1 0 1592 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1522732896
transform 1 0 1608 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_2
timestamp 1522732896
transform 1 0 1624 0 1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_29
timestamp 1522732896
transform 1 0 1640 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_94
timestamp 1522732896
transform 1 0 1704 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_318
timestamp 1522732896
transform -1 0 1832 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_29
timestamp 1522732896
transform 1 0 1832 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_319
timestamp 1522732896
transform 1 0 1896 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_19
timestamp 1522732896
transform -1 0 2024 0 1 3410
box 0 0 64 200
use INVX1  INVX1_26
timestamp 1522732896
transform 1 0 2024 0 1 3410
box 0 0 32 200
use AOI21X1  AOI21X1_20
timestamp 1522732896
transform 1 0 2056 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_360
timestamp 1522732896
transform -1 0 2184 0 1 3410
box 0 0 64 200
use INVX1  INVX1_21
timestamp 1522732896
transform -1 0 2216 0 1 3410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_102
timestamp 1522732896
transform -1 0 2408 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_348
timestamp 1522732896
transform 1 0 2408 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_19
timestamp 1522732896
transform -1 0 2536 0 1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_11
timestamp 1522732896
transform 1 0 2536 0 1 3410
box 0 0 80 200
use OAI22X1  OAI22X1_22
timestamp 1522732896
transform 1 0 2616 0 1 3410
box 0 0 80 200
use INVX2  INVX2_16
timestamp 1522732896
transform -1 0 2728 0 1 3410
box 0 0 32 200
use AOI21X1  AOI21X1_54
timestamp 1522732896
transform -1 0 2792 0 1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_21
timestamp 1522732896
transform 1 0 2792 0 1 3410
box 0 0 80 200
use OAI22X1  OAI22X1_12
timestamp 1522732896
transform 1 0 2872 0 1 3410
box 0 0 80 200
use OAI22X1  OAI22X1_23
timestamp 1522732896
transform 1 0 2952 0 1 3410
box 0 0 80 200
use OAI22X1  OAI22X1_14
timestamp 1522732896
transform 1 0 3032 0 1 3410
box 0 0 80 200
use FILL  FILL_17_1_0
timestamp 1522732896
transform -1 0 3128 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1522732896
transform -1 0 3144 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_2
timestamp 1522732896
transform -1 0 3160 0 1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_55
timestamp 1522732896
transform -1 0 3224 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_53
timestamp 1522732896
transform -1 0 3288 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_154
timestamp 1522732896
transform -1 0 3352 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_31
timestamp 1522732896
transform -1 0 3416 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_93
timestamp 1522732896
transform -1 0 3480 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_28
timestamp 1522732896
transform -1 0 3544 0 1 3410
box 0 0 64 200
use INVX4  INVX4_5
timestamp 1522732896
transform 1 0 3544 0 1 3410
box 0 0 48 200
use OAI22X1  OAI22X1_13
timestamp 1522732896
transform 1 0 3592 0 1 3410
box 0 0 80 200
use NAND3X1  NAND3X1_116
timestamp 1522732896
transform -1 0 3736 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_104
timestamp 1522732896
transform 1 0 3736 0 1 3410
box 0 0 64 200
use BUFX2  BUFX2_5
timestamp 1522732896
transform 1 0 3800 0 1 3410
box 0 0 48 200
use MUX2X1  MUX2X1_12
timestamp 1522732896
transform -1 0 3944 0 1 3410
box 0 0 96 200
use NAND3X1  NAND3X1_103
timestamp 1522732896
transform 1 0 3944 0 1 3410
box 0 0 64 200
use INVX1  INVX1_75
timestamp 1522732896
transform -1 0 4040 0 1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_115
timestamp 1522732896
transform -1 0 4104 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_118
timestamp 1522732896
transform 1 0 4104 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_135
timestamp 1522732896
transform -1 0 4216 0 1 3410
box 0 0 48 200
use MUX2X1  MUX2X1_16
timestamp 1522732896
transform 1 0 4216 0 1 3410
box 0 0 96 200
use INVX1  INVX1_87
timestamp 1522732896
transform -1 0 4344 0 1 3410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1522732896
transform -1 0 4536 0 1 3410
box 0 0 192 200
use INVX1  INVX1_70
timestamp 1522732896
transform -1 0 4568 0 1 3410
box 0 0 32 200
use MUX2X1  MUX2X1_11
timestamp 1522732896
transform 1 0 4568 0 1 3410
box 0 0 96 200
use FILL  FILL_17_2_0
timestamp 1522732896
transform -1 0 4680 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1522732896
transform -1 0 4696 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_2
timestamp 1522732896
transform -1 0 4712 0 1 3410
box 0 0 16 200
use INVX1  INVX1_78
timestamp 1522732896
transform -1 0 4744 0 1 3410
box 0 0 32 200
use INVX1  INVX1_90
timestamp 1522732896
transform -1 0 4776 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_284
timestamp 1522732896
transform 1 0 4776 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_182
timestamp 1522732896
transform -1 0 4888 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1522732896
transform -1 0 5080 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_224
timestamp 1522732896
transform 1 0 5080 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_422
timestamp 1522732896
transform 1 0 5128 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_423
timestamp 1522732896
transform -1 0 5256 0 1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_57
timestamp 1522732896
transform 1 0 5256 0 1 3410
box 0 0 80 200
use INVX1  INVX1_180
timestamp 1522732896
transform 1 0 5336 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_235
timestamp 1522732896
transform -1 0 5416 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_52
timestamp 1522732896
transform -1 0 5496 0 1 3410
box 0 0 80 200
use AND2X2  AND2X2_48
timestamp 1522732896
transform -1 0 5560 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_402
timestamp 1522732896
transform 1 0 5560 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_401
timestamp 1522732896
transform -1 0 5688 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_232
timestamp 1522732896
transform -1 0 5736 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_405
timestamp 1522732896
transform 1 0 5736 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_404
timestamp 1522732896
transform -1 0 5864 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_166
timestamp 1522732896
transform 1 0 5864 0 1 3410
box 0 0 64 200
use INVX1  INVX1_176
timestamp 1522732896
transform 1 0 5928 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_411
timestamp 1522732896
transform 1 0 5960 0 1 3410
box 0 0 64 200
use INVX1  INVX1_175
timestamp 1522732896
transform -1 0 6056 0 1 3410
box 0 0 32 200
use INVX1  INVX1_170
timestamp 1522732896
transform -1 0 6088 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_229
timestamp 1522732896
transform -1 0 6136 0 1 3410
box 0 0 48 200
use INVX1  INVX1_163
timestamp 1522732896
transform -1 0 6168 0 1 3410
box 0 0 32 200
use INVX1  INVX1_178
timestamp 1522732896
transform -1 0 6200 0 1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_218
timestamp 1522732896
transform -1 0 6248 0 1 3410
box 0 0 48 200
use FILL  FILL_18_1
timestamp 1522732896
transform 1 0 6248 0 1 3410
box 0 0 16 200
use FILL  FILL_18_2
timestamp 1522732896
transform 1 0 6264 0 1 3410
box 0 0 16 200
use FILL  FILL_18_3
timestamp 1522732896
transform 1 0 6280 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_113
timestamp 1522732896
transform 1 0 8 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_210
timestamp 1522732896
transform 1 0 200 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_118
timestamp 1522732896
transform 1 0 248 0 -1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_10
timestamp 1522732896
transform -1 0 504 0 -1 3410
box 0 0 64 200
use INVX2  INVX2_13
timestamp 1522732896
transform 1 0 504 0 -1 3410
box 0 0 32 200
use INVX2  INVX2_14
timestamp 1522732896
transform 1 0 536 0 -1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_21
timestamp 1522732896
transform -1 0 632 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_17
timestamp 1522732896
transform 1 0 632 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_26
timestamp 1522732896
transform 1 0 680 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_22
timestamp 1522732896
transform -1 0 792 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_5
timestamp 1522732896
transform -1 0 856 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_14
timestamp 1522732896
transform -1 0 920 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_25
timestamp 1522732896
transform -1 0 984 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_35
timestamp 1522732896
transform -1 0 1048 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_11
timestamp 1522732896
transform 1 0 1048 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_5
timestamp 1522732896
transform -1 0 1176 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_10
timestamp 1522732896
transform 1 0 1176 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_18
timestamp 1522732896
transform 1 0 1240 0 -1 3410
box 0 0 48 200
use AOI21X1  AOI21X1_28
timestamp 1522732896
transform 1 0 1288 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_35
timestamp 1522732896
transform -1 0 1416 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_32
timestamp 1522732896
transform -1 0 1464 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_29
timestamp 1522732896
transform 1 0 1464 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_30
timestamp 1522732896
transform -1 0 1576 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_0_0
timestamp 1522732896
transform 1 0 1576 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1522732896
transform 1 0 1592 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_2
timestamp 1522732896
transform 1 0 1608 0 -1 3410
box 0 0 16 200
use NOR2X1  NOR2X1_33
timestamp 1522732896
transform 1 0 1624 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_47
timestamp 1522732896
transform 1 0 1672 0 -1 3410
box 0 0 80 200
use BUFX4  BUFX4_34
timestamp 1522732896
transform 1 0 1752 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_44
timestamp 1522732896
transform 1 0 1816 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_317
timestamp 1522732896
transform -1 0 1960 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_32
timestamp 1522732896
transform 1 0 1960 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_349
timestamp 1522732896
transform -1 0 2088 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_350
timestamp 1522732896
transform -1 0 2152 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_108
timestamp 1522732896
transform -1 0 2216 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_353
timestamp 1522732896
transform -1 0 2280 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_357
timestamp 1522732896
transform 1 0 2280 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_109
timestamp 1522732896
transform 1 0 2344 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_110
timestamp 1522732896
transform 1 0 2408 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_197
timestamp 1522732896
transform -1 0 2520 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_347
timestamp 1522732896
transform 1 0 2520 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_214
timestamp 1522732896
transform -1 0 2632 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_358
timestamp 1522732896
transform -1 0 2696 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_354
timestamp 1522732896
transform -1 0 2760 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_137
timestamp 1522732896
transform 1 0 2760 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_141
timestamp 1522732896
transform -1 0 2872 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_138
timestamp 1522732896
transform 1 0 2872 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_153
timestamp 1522732896
transform -1 0 2984 0 -1 3410
box 0 0 64 200
use INVX2  INVX2_41
timestamp 1522732896
transform -1 0 3016 0 -1 3410
box 0 0 32 200
use OAI22X1  OAI22X1_15
timestamp 1522732896
transform 1 0 3016 0 -1 3410
box 0 0 80 200
use INVX1  INVX1_123
timestamp 1522732896
transform 1 0 3096 0 -1 3410
box 0 0 32 200
use FILL  FILL_16_1_0
timestamp 1522732896
transform 1 0 3128 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1522732896
transform 1 0 3144 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_2
timestamp 1522732896
transform 1 0 3160 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_31
timestamp 1522732896
transform 1 0 3176 0 -1 3410
box 0 0 64 200
use INVX2  INVX2_35
timestamp 1522732896
transform -1 0 3272 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_176
timestamp 1522732896
transform -1 0 3336 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_157
timestamp 1522732896
transform 1 0 3336 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_171
timestamp 1522732896
transform 1 0 3400 0 -1 3410
box 0 0 64 200
use BUFX2  BUFX2_34
timestamp 1522732896
transform 1 0 3464 0 -1 3410
box 0 0 48 200
use INVX2  INVX2_21
timestamp 1522732896
transform -1 0 3544 0 -1 3410
box 0 0 32 200
use AOI22X1  AOI22X1_31
timestamp 1522732896
transform 1 0 3544 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_192
timestamp 1522732896
transform 1 0 3624 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_146
timestamp 1522732896
transform 1 0 3688 0 -1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_156
timestamp 1522732896
transform 1 0 3736 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_30
timestamp 1522732896
transform -1 0 3864 0 -1 3410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1522732896
transform 1 0 3864 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_128
timestamp 1522732896
transform -1 0 4104 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_134
timestamp 1522732896
transform -1 0 4152 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_133
timestamp 1522732896
transform -1 0 4200 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_88
timestamp 1522732896
transform -1 0 4232 0 -1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_171
timestamp 1522732896
transform 1 0 4232 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_239
timestamp 1522732896
transform -1 0 4344 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1522732896
transform -1 0 4536 0 -1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1522732896
transform -1 0 4728 0 -1 3410
box 0 0 192 200
use FILL  FILL_16_2_0
timestamp 1522732896
transform 1 0 4728 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1522732896
transform 1 0 4744 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_2
timestamp 1522732896
transform 1 0 4760 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_287
timestamp 1522732896
transform 1 0 4776 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_185
timestamp 1522732896
transform -1 0 4888 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1522732896
transform -1 0 5080 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_245
timestamp 1522732896
transform 1 0 5080 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_464
timestamp 1522732896
transform -1 0 5192 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_223
timestamp 1522732896
transform -1 0 5240 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_214
timestamp 1522732896
transform 1 0 5240 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_400
timestamp 1522732896
transform 1 0 5288 0 -1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_55
timestamp 1522732896
transform -1 0 5432 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_436
timestamp 1522732896
transform 1 0 5432 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_435
timestamp 1522732896
transform -1 0 5560 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_403
timestamp 1522732896
transform -1 0 5624 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_171
timestamp 1522732896
transform 1 0 5624 0 -1 3410
box 0 0 32 200
use INVX1  INVX1_200
timestamp 1522732896
transform 1 0 5656 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_452
timestamp 1522732896
transform 1 0 5688 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_240
timestamp 1522732896
transform -1 0 5800 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_239
timestamp 1522732896
transform -1 0 5848 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_185
timestamp 1522732896
transform 1 0 5848 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_457
timestamp 1522732896
transform 1 0 5880 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_126
timestamp 1522732896
transform 1 0 5944 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_453
timestamp 1522732896
transform 1 0 6008 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_174
timestamp 1522732896
transform 1 0 6072 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_61
timestamp 1522732896
transform -1 0 6216 0 -1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_234
timestamp 1522732896
transform -1 0 6264 0 -1 3410
box 0 0 48 200
use FILL  FILL_17_1
timestamp 1522732896
transform -1 0 6280 0 -1 3410
box 0 0 16 200
use FILL  FILL_17_2
timestamp 1522732896
transform -1 0 6296 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_112
timestamp 1522732896
transform 1 0 8 0 1 3010
box 0 0 192 200
use OAI22X1  OAI22X1_47
timestamp 1522732896
transform 1 0 200 0 1 3010
box 0 0 80 200
use NOR2X1  NOR2X1_217
timestamp 1522732896
transform 1 0 280 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_25
timestamp 1522732896
transform 1 0 328 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_162
timestamp 1522732896
transform 1 0 392 0 1 3010
box 0 0 64 200
use INVX1  INVX1_158
timestamp 1522732896
transform -1 0 488 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_35
timestamp 1522732896
transform -1 0 536 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_23
timestamp 1522732896
transform -1 0 600 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_376
timestamp 1522732896
transform 1 0 600 0 1 3010
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1522732896
transform -1 0 696 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_8
timestamp 1522732896
transform -1 0 776 0 1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_36
timestamp 1522732896
transform -1 0 840 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_27
timestamp 1522732896
transform 1 0 840 0 1 3010
box 0 0 48 200
use AND2X2  AND2X2_6
timestamp 1522732896
transform -1 0 952 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_24
timestamp 1522732896
transform 1 0 952 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_18
timestamp 1522732896
transform -1 0 1080 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_7
timestamp 1522732896
transform -1 0 1160 0 1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_27
timestamp 1522732896
transform 1 0 1160 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_32
timestamp 1522732896
transform 1 0 1224 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_95
timestamp 1522732896
transform 1 0 1288 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_20
timestamp 1522732896
transform 1 0 1480 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_25
timestamp 1522732896
transform 1 0 1528 0 1 3010
box 0 0 48 200
use FILL  FILL_15_0_0
timestamp 1522732896
transform 1 0 1576 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1522732896
transform 1 0 1592 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_2
timestamp 1522732896
transform 1 0 1608 0 1 3010
box 0 0 16 200
use OAI21X1  OAI21X1_21
timestamp 1522732896
transform 1 0 1624 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_24
timestamp 1522732896
transform -1 0 1736 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_341
timestamp 1522732896
transform 1 0 1736 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_342
timestamp 1522732896
transform -1 0 1864 0 1 3010
box 0 0 64 200
use INVX1  INVX1_155
timestamp 1522732896
transform 1 0 1864 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_320
timestamp 1522732896
transform -1 0 1960 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_11
timestamp 1522732896
transform 1 0 1960 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_337
timestamp 1522732896
transform 1 0 2024 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_200
timestamp 1522732896
transform -1 0 2136 0 1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_104
timestamp 1522732896
transform -1 0 2200 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_199
timestamp 1522732896
transform -1 0 2248 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_194
timestamp 1522732896
transform 1 0 2248 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_338
timestamp 1522732896
transform -1 0 2360 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_201
timestamp 1522732896
transform -1 0 2408 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_361
timestamp 1522732896
transform 1 0 2408 0 1 3010
box 0 0 64 200
use OAI22X1  OAI22X1_30
timestamp 1522732896
transform 1 0 2472 0 1 3010
box 0 0 80 200
use OAI22X1  OAI22X1_29
timestamp 1522732896
transform 1 0 2552 0 1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_159
timestamp 1522732896
transform -1 0 2696 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_345
timestamp 1522732896
transform -1 0 2760 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_107
timestamp 1522732896
transform 1 0 2760 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_198
timestamp 1522732896
transform -1 0 2888 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1522732896
transform 1 0 2888 0 1 3010
box 0 0 192 200
use AND2X2  AND2X2_38
timestamp 1522732896
transform -1 0 3144 0 1 3010
box 0 0 64 200
use FILL  FILL_15_1_0
timestamp 1522732896
transform -1 0 3160 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1522732896
transform -1 0 3176 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_2
timestamp 1522732896
transform -1 0 3192 0 1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_64
timestamp 1522732896
transform -1 0 3256 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_159
timestamp 1522732896
transform 1 0 3256 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_158
timestamp 1522732896
transform 1 0 3320 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1522732896
transform -1 0 3448 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_73
timestamp 1522732896
transform -1 0 3640 0 1 3010
box 0 0 192 200
use INVX2  INVX2_11
timestamp 1522732896
transform 1 0 3640 0 1 3010
box 0 0 32 200
use INVX1  INVX1_122
timestamp 1522732896
transform -1 0 3704 0 1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_73
timestamp 1522732896
transform -1 0 3768 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_155
timestamp 1522732896
transform 1 0 3768 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_147
timestamp 1522732896
transform -1 0 3864 0 1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_32
timestamp 1522732896
transform -1 0 3944 0 1 3010
box 0 0 80 200
use XNOR2X1  XNOR2X1_2
timestamp 1522732896
transform -1 0 4056 0 1 3010
box 0 0 112 200
use OAI21X1  OAI21X1_193
timestamp 1522732896
transform 1 0 4056 0 1 3010
box 0 0 64 200
use BUFX2  BUFX2_4
timestamp 1522732896
transform -1 0 4168 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_150
timestamp 1522732896
transform -1 0 4232 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_16
timestamp 1522732896
transform -1 0 4296 0 1 3010
box 0 0 64 200
use INVX1  INVX1_121
timestamp 1522732896
transform -1 0 4328 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_286
timestamp 1522732896
transform 1 0 4328 0 1 3010
box 0 0 64 200
use INVX1  INVX1_86
timestamp 1522732896
transform -1 0 4424 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_184
timestamp 1522732896
transform -1 0 4472 0 1 3010
box 0 0 48 200
use INVX1  INVX1_165
timestamp 1522732896
transform 1 0 4472 0 1 3010
box 0 0 32 200
use INVX1  INVX1_76
timestamp 1522732896
transform -1 0 4536 0 1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1522732896
transform -1 0 4728 0 1 3010
box 0 0 192 200
use FILL  FILL_15_2_0
timestamp 1522732896
transform 1 0 4728 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1522732896
transform 1 0 4744 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_2
timestamp 1522732896
transform 1 0 4760 0 1 3010
box 0 0 16 200
use OAI21X1  OAI21X1_236
timestamp 1522732896
transform 1 0 4776 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_168
timestamp 1522732896
transform -1 0 4888 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_130
timestamp 1522732896
transform -1 0 5080 0 1 3010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_134
timestamp 1522732896
transform -1 0 5272 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_469
timestamp 1522732896
transform -1 0 5336 0 1 3010
box 0 0 64 200
use INVX1  INVX1_164
timestamp 1522732896
transform 1 0 5336 0 1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_230
timestamp 1522732896
transform -1 0 5416 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_396
timestamp 1522732896
transform -1 0 5480 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_51
timestamp 1522732896
transform -1 0 5560 0 1 3010
box 0 0 80 200
use INVX1  INVX1_194
timestamp 1522732896
transform 1 0 5560 0 1 3010
box 0 0 32 200
use INVX1  INVX1_193
timestamp 1522732896
transform 1 0 5592 0 1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_128
timestamp 1522732896
transform 1 0 5624 0 1 3010
box 0 0 64 200
use INVX1  INVX1_169
timestamp 1522732896
transform 1 0 5688 0 1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_130
timestamp 1522732896
transform -1 0 5784 0 1 3010
box 0 0 64 200
use INVX1  INVX1_167
timestamp 1522732896
transform 1 0 5784 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_437
timestamp 1522732896
transform 1 0 5816 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_399
timestamp 1522732896
transform -1 0 5944 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_231
timestamp 1522732896
transform -1 0 5992 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_237
timestamp 1522732896
transform -1 0 6040 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_241
timestamp 1522732896
transform -1 0 6088 0 1 3010
box 0 0 48 200
use INVX1  INVX1_199
timestamp 1522732896
transform -1 0 6120 0 1 3010
box 0 0 32 200
use INVX1  INVX1_196
timestamp 1522732896
transform 1 0 6120 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_449
timestamp 1522732896
transform -1 0 6216 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_447
timestamp 1522732896
transform 1 0 6216 0 1 3010
box 0 0 64 200
use FILL  FILL_16_1
timestamp 1522732896
transform 1 0 6280 0 1 3010
box 0 0 16 200
use OAI22X1  OAI22X1_48
timestamp 1522732896
transform 1 0 8 0 -1 3010
box 0 0 80 200
use AND2X2  AND2X2_46
timestamp 1522732896
transform -1 0 152 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_377
timestamp 1522732896
transform -1 0 216 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_208
timestamp 1522732896
transform 1 0 216 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_160
timestamp 1522732896
transform -1 0 328 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_19
timestamp 1522732896
transform 1 0 328 0 -1 3010
box 0 0 48 200
use AND2X2  AND2X2_4
timestamp 1522732896
transform 1 0 376 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1522732896
transform 1 0 440 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_36
timestamp 1522732896
transform -1 0 552 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_28
timestamp 1522732896
transform 1 0 552 0 -1 3010
box 0 0 32 200
use OAI22X1  OAI22X1_4
timestamp 1522732896
transform -1 0 664 0 -1 3010
box 0 0 80 200
use NOR2X1  NOR2X1_218
timestamp 1522732896
transform -1 0 712 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_378
timestamp 1522732896
transform -1 0 776 0 -1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_16
timestamp 1522732896
transform -1 0 840 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_35
timestamp 1522732896
transform -1 0 904 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_37
timestamp 1522732896
transform -1 0 968 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_36
timestamp 1522732896
transform 1 0 968 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_28
timestamp 1522732896
transform -1 0 1080 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_18
timestamp 1522732896
transform 1 0 1080 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_7
timestamp 1522732896
transform -1 0 1176 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_75
timestamp 1522732896
transform 1 0 1176 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1522732896
transform 1 0 1240 0 -1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_8
timestamp 1522732896
transform -1 0 1368 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_38
timestamp 1522732896
transform -1 0 1432 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_39
timestamp 1522732896
transform 1 0 1432 0 -1 3010
box 0 0 64 200
use BUFX2  BUFX2_11
timestamp 1522732896
transform -1 0 1544 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_34
timestamp 1522732896
transform 1 0 1544 0 -1 3010
box 0 0 48 200
use FILL  FILL_14_0_0
timestamp 1522732896
transform -1 0 1608 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1522732896
transform -1 0 1624 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_2
timestamp 1522732896
transform -1 0 1640 0 -1 3010
box 0 0 16 200
use AOI22X1  AOI22X1_50
timestamp 1522732896
transform -1 0 1720 0 -1 3010
box 0 0 80 200
use AOI21X1  AOI21X1_106
timestamp 1522732896
transform 1 0 1720 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_49
timestamp 1522732896
transform 1 0 1784 0 -1 3010
box 0 0 80 200
use OR2X2  OR2X2_25
timestamp 1522732896
transform -1 0 1928 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_23
timestamp 1522732896
transform 1 0 1928 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_364
timestamp 1522732896
transform 1 0 1992 0 -1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_112
timestamp 1522732896
transform -1 0 2120 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_54
timestamp 1522732896
transform 1 0 2120 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_24
timestamp 1522732896
transform -1 0 2248 0 -1 3010
box 0 0 64 200
use OAI22X1  OAI22X1_32
timestamp 1522732896
transform -1 0 2328 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_362
timestamp 1522732896
transform 1 0 2328 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_106
timestamp 1522732896
transform 1 0 2392 0 -1 3010
box 0 0 192 200
use AOI21X1  AOI21X1_111
timestamp 1522732896
transform -1 0 2648 0 -1 3010
box 0 0 64 200
use INVX2  INVX2_22
timestamp 1522732896
transform 1 0 2648 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_16
timestamp 1522732896
transform -1 0 2728 0 -1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_63
timestamp 1522732896
transform -1 0 2792 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_37
timestamp 1522732896
transform 1 0 2792 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_143
timestamp 1522732896
transform 1 0 2856 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_148
timestamp 1522732896
transform 1 0 2904 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_9
timestamp 1522732896
transform 1 0 2952 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_67
timestamp 1522732896
transform -1 0 3048 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_160
timestamp 1522732896
transform -1 0 3112 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_1_0
timestamp 1522732896
transform 1 0 3112 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1522732896
transform 1 0 3128 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_2
timestamp 1522732896
transform 1 0 3144 0 -1 3010
box 0 0 16 200
use OAI22X1  OAI22X1_24
timestamp 1522732896
transform 1 0 3160 0 -1 3010
box 0 0 80 200
use AOI21X1  AOI21X1_56
timestamp 1522732896
transform -1 0 3304 0 -1 3010
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1522732896
transform 1 0 3304 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_57
timestamp 1522732896
transform 1 0 3336 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_191
timestamp 1522732896
transform -1 0 3464 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_195
timestamp 1522732896
transform -1 0 3528 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_33
timestamp 1522732896
transform 1 0 3528 0 -1 3010
box 0 0 80 200
use AOI21X1  AOI21X1_74
timestamp 1522732896
transform -1 0 3672 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_150
timestamp 1522732896
transform 1 0 3672 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_127
timestamp 1522732896
transform 1 0 3720 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_196
timestamp 1522732896
transform -1 0 3816 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_149
timestamp 1522732896
transform 1 0 3816 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_157
timestamp 1522732896
transform 1 0 3864 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_158
timestamp 1522732896
transform 1 0 3912 0 -1 3010
box 0 0 48 200
use MUX2X1  MUX2X1_14
timestamp 1522732896
transform 1 0 3960 0 -1 3010
box 0 0 96 200
use XNOR2X1  XNOR2X1_4
timestamp 1522732896
transform 1 0 4056 0 -1 3010
box 0 0 112 200
use XNOR2X1  XNOR2X1_3
timestamp 1522732896
transform -1 0 4280 0 -1 3010
box 0 0 112 200
use NAND2X1  NAND2X1_145
timestamp 1522732896
transform 1 0 4280 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1522732896
transform 1 0 4328 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_144
timestamp 1522732896
transform 1 0 4520 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_154
timestamp 1522732896
transform -1 0 4616 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_132
timestamp 1522732896
transform 1 0 4616 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_2_0
timestamp 1522732896
transform 1 0 4680 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1522732896
transform 1 0 4696 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_2
timestamp 1522732896
transform 1 0 4712 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_20
timestamp 1522732896
transform 1 0 4728 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_128
timestamp 1522732896
transform 1 0 4792 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_243
timestamp 1522732896
transform 1 0 4984 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_460
timestamp 1522732896
transform -1 0 5096 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_66
timestamp 1522732896
transform -1 0 5160 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_249
timestamp 1522732896
transform 1 0 5160 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_398
timestamp 1522732896
transform 1 0 5208 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_395
timestamp 1522732896
transform 1 0 5272 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_166
timestamp 1522732896
transform 1 0 5336 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_121
timestamp 1522732896
transform 1 0 5368 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_238
timestamp 1522732896
transform 1 0 5432 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_192
timestamp 1522732896
transform -1 0 5512 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_444
timestamp 1522732896
transform 1 0 5512 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_443
timestamp 1522732896
transform -1 0 5640 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_59
timestamp 1522732896
transform -1 0 5720 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_446
timestamp 1522732896
transform 1 0 5720 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_169
timestamp 1522732896
transform 1 0 5784 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_170
timestamp 1522732896
transform -1 0 5912 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_39
timestamp 1522732896
transform -1 0 5976 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_450
timestamp 1522732896
transform 1 0 5976 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_230
timestamp 1522732896
transform 1 0 6040 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_173
timestamp 1522732896
transform -1 0 6152 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_454
timestamp 1522732896
transform 1 0 6152 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_198
timestamp 1522732896
transform -1 0 6248 0 -1 3010
box 0 0 32 200
use INVX1  INVX1_197
timestamp 1522732896
transform 1 0 6248 0 -1 3010
box 0 0 32 200
use FILL  FILL_15_1
timestamp 1522732896
transform -1 0 6296 0 -1 3010
box 0 0 16 200
use NOR3X1  NOR3X1_15
timestamp 1522732896
transform -1 0 136 0 1 2610
box 0 0 128 200
use NOR2X1  NOR2X1_219
timestamp 1522732896
transform 1 0 136 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_379
timestamp 1522732896
transform -1 0 248 0 1 2610
box 0 0 64 200
use INVX1  INVX1_159
timestamp 1522732896
transform -1 0 280 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_381
timestamp 1522732896
transform -1 0 344 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_3
timestamp 1522732896
transform 1 0 344 0 1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_7
timestamp 1522732896
transform -1 0 488 0 1 2610
box 0 0 64 200
use INVX2  INVX2_4
timestamp 1522732896
transform 1 0 488 0 1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_207
timestamp 1522732896
transform 1 0 520 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_216
timestamp 1522732896
transform -1 0 616 0 1 2610
box 0 0 48 200
use OAI22X1  OAI22X1_46
timestamp 1522732896
transform -1 0 696 0 1 2610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_111
timestamp 1522732896
transform 1 0 696 0 1 2610
box 0 0 192 200
use INVX2  INVX2_12
timestamp 1522732896
transform -1 0 920 0 1 2610
box 0 0 32 200
use NAND3X1  NAND3X1_19
timestamp 1522732896
transform -1 0 984 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_27
timestamp 1522732896
transform -1 0 1064 0 1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_20
timestamp 1522732896
transform -1 0 1128 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_20
timestamp 1522732896
transform 1 0 1128 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1522732896
transform -1 0 1256 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_4
timestamp 1522732896
transform -1 0 1320 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_3
timestamp 1522732896
transform -1 0 1384 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_2
timestamp 1522732896
transform 1 0 1384 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_32
timestamp 1522732896
transform 1 0 1448 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1522732896
transform -1 0 1560 0 1 2610
box 0 0 48 200
use FILL  FILL_13_0_0
timestamp 1522732896
transform -1 0 1576 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1522732896
transform -1 0 1592 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_2
timestamp 1522732896
transform -1 0 1608 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_33
timestamp 1522732896
transform -1 0 1672 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_31
timestamp 1522732896
transform 1 0 1672 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_32
timestamp 1522732896
transform -1 0 1800 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1522732896
transform 1 0 1800 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_1
timestamp 1522732896
transform -1 0 1928 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_33
timestamp 1522732896
transform 1 0 1928 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_363
timestamp 1522732896
transform 1 0 1992 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_365
timestamp 1522732896
transform 1 0 2056 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_371
timestamp 1522732896
transform 1 0 2120 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_204
timestamp 1522732896
transform 1 0 2184 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_369
timestamp 1522732896
transform 1 0 2232 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_203
timestamp 1522732896
transform 1 0 2296 0 1 2610
box 0 0 48 200
use INVX2  INVX2_44
timestamp 1522732896
transform 1 0 2344 0 1 2610
box 0 0 32 200
use AOI21X1  AOI21X1_113
timestamp 1522732896
transform 1 0 2376 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_368
timestamp 1522732896
transform -1 0 2504 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_202
timestamp 1522732896
transform 1 0 2504 0 1 2610
box 0 0 48 200
use OAI22X1  OAI22X1_43
timestamp 1522732896
transform 1 0 2552 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_366
timestamp 1522732896
transform -1 0 2696 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_107
timestamp 1522732896
transform 1 0 2696 0 1 2610
box 0 0 192 200
use INVX1  INVX1_91
timestamp 1522732896
transform 1 0 2888 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_175
timestamp 1522732896
transform -1 0 2984 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1522732896
transform 1 0 2984 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_7
timestamp 1522732896
transform 1 0 3048 0 1 2610
box 0 0 48 200
use FILL  FILL_13_1_0
timestamp 1522732896
transform 1 0 3096 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1522732896
transform 1 0 3112 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_2
timestamp 1522732896
transform 1 0 3128 0 1 2610
box 0 0 16 200
use INVX8  INVX8_3
timestamp 1522732896
transform 1 0 3144 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_5
timestamp 1522732896
transform -1 0 3288 0 1 2610
box 0 0 64 200
use INVX1  INVX1_113
timestamp 1522732896
transform 1 0 3288 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_170
timestamp 1522732896
transform -1 0 3384 0 1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_25
timestamp 1522732896
transform 1 0 3384 0 1 2610
box 0 0 80 200
use INVX2  INVX2_23
timestamp 1522732896
transform -1 0 3496 0 1 2610
box 0 0 32 200
use INVX1  INVX1_128
timestamp 1522732896
transform 1 0 3496 0 1 2610
box 0 0 32 200
use OAI22X1  OAI22X1_16
timestamp 1522732896
transform 1 0 3528 0 1 2610
box 0 0 80 200
use OAI22X1  OAI22X1_17
timestamp 1522732896
transform 1 0 3608 0 1 2610
box 0 0 80 200
use MUX2X1  MUX2X1_19
timestamp 1522732896
transform 1 0 3688 0 1 2610
box 0 0 96 200
use OAI21X1  OAI21X1_197
timestamp 1522732896
transform -1 0 3848 0 1 2610
box 0 0 64 200
use INVX1  INVX1_66
timestamp 1522732896
transform -1 0 3880 0 1 2610
box 0 0 32 200
use INVX1  INVX1_126
timestamp 1522732896
transform 1 0 3880 0 1 2610
box 0 0 32 200
use XNOR2X1  XNOR2X1_7
timestamp 1522732896
transform -1 0 4024 0 1 2610
box 0 0 112 200
use NOR2X1  NOR2X1_226
timestamp 1522732896
transform -1 0 4072 0 1 2610
box 0 0 48 200
use OR2X2  OR2X2_38
timestamp 1522732896
transform -1 0 4136 0 1 2610
box 0 0 64 200
use XNOR2X1  XNOR2X1_5
timestamp 1522732896
transform -1 0 4248 0 1 2610
box 0 0 112 200
use INVX2  INVX2_26
timestamp 1522732896
transform -1 0 4280 0 1 2610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_78
timestamp 1522732896
transform -1 0 4472 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_274
timestamp 1522732896
transform 1 0 4472 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_80
timestamp 1522732896
transform 1 0 4536 0 1 2610
box 0 0 192 200
use FILL  FILL_13_2_0
timestamp 1522732896
transform 1 0 4728 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1522732896
transform 1 0 4744 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_2
timestamp 1522732896
transform 1 0 4760 0 1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_23
timestamp 1522732896
transform 1 0 4776 0 1 2610
box 0 0 96 200
use INVX1  INVX1_146
timestamp 1522732896
transform -1 0 4904 0 1 2610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_82
timestamp 1522732896
transform -1 0 5096 0 1 2610
box 0 0 192 200
use MUX2X1  MUX2X1_22
timestamp 1522732896
transform 1 0 5096 0 1 2610
box 0 0 96 200
use INVX1  INVX1_145
timestamp 1522732896
transform -1 0 5224 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_397
timestamp 1522732896
transform 1 0 5224 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_81
timestamp 1522732896
transform 1 0 5288 0 1 2610
box 0 0 192 200
use NOR2X1  NOR2X1_237
timestamp 1522732896
transform 1 0 5480 0 1 2610
box 0 0 48 200
use INVX1  INVX1_186
timestamp 1522732896
transform -1 0 5560 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_439
timestamp 1522732896
transform 1 0 5560 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_438
timestamp 1522732896
transform -1 0 5688 0 1 2610
box 0 0 64 200
use INVX1  INVX1_187
timestamp 1522732896
transform 1 0 5688 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_445
timestamp 1522732896
transform -1 0 5784 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_63
timestamp 1522732896
transform 1 0 5784 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_440
timestamp 1522732896
transform 1 0 5864 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_441
timestamp 1522732896
transform 1 0 5928 0 1 2610
box 0 0 64 200
use INVX4  INVX4_8
timestamp 1522732896
transform -1 0 6040 0 1 2610
box 0 0 48 200
use INVX1  INVX1_190
timestamp 1522732896
transform 1 0 6040 0 1 2610
box 0 0 32 200
use AOI21X1  AOI21X1_132
timestamp 1522732896
transform -1 0 6136 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_238
timestamp 1522732896
transform 1 0 6136 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_448
timestamp 1522732896
transform 1 0 6184 0 1 2610
box 0 0 64 200
use FILL  FILL_14_1
timestamp 1522732896
transform 1 0 6248 0 1 2610
box 0 0 16 200
use FILL  FILL_14_2
timestamp 1522732896
transform 1 0 6264 0 1 2610
box 0 0 16 200
use FILL  FILL_14_3
timestamp 1522732896
transform 1 0 6280 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_3
timestamp 1522732896
transform 1 0 8 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_36
timestamp 1522732896
transform 1 0 72 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_115
timestamp 1522732896
transform -1 0 200 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_116
timestamp 1522732896
transform 1 0 200 0 -1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_49
timestamp 1522732896
transform -1 0 344 0 -1 2610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_115
timestamp 1522732896
transform 1 0 344 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_6
timestamp 1522732896
transform -1 0 584 0 -1 2610
box 0 0 48 200
use AND2X2  AND2X2_8
timestamp 1522732896
transform -1 0 648 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1522732896
transform 1 0 648 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_34
timestamp 1522732896
transform 1 0 712 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_36
timestamp 1522732896
transform 1 0 776 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_13
timestamp 1522732896
transform -1 0 920 0 -1 2610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_125
timestamp 1522732896
transform 1 0 920 0 -1 2610
box 0 0 192 200
use INVX1  INVX1_30
timestamp 1522732896
transform 1 0 1112 0 -1 2610
box 0 0 32 200
use AOI22X1  AOI22X1_2
timestamp 1522732896
transform 1 0 1144 0 -1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_25
timestamp 1522732896
transform 1 0 1224 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_26
timestamp 1522732896
transform 1 0 1272 0 -1 2610
box 0 0 48 200
use OAI22X1  OAI22X1_3
timestamp 1522732896
transform -1 0 1400 0 -1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_6
timestamp 1522732896
transform -1 0 1464 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_39
timestamp 1522732896
transform -1 0 1528 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_34
timestamp 1522732896
transform 1 0 1528 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_0_0
timestamp 1522732896
transform -1 0 1608 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1522732896
transform -1 0 1624 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_2
timestamp 1522732896
transform -1 0 1640 0 -1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_39
timestamp 1522732896
transform -1 0 1704 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_11
timestamp 1522732896
transform -1 0 1784 0 -1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_35
timestamp 1522732896
transform 1 0 1784 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_8
timestamp 1522732896
transform -1 0 1880 0 -1 2610
box 0 0 48 200
use AOI21X1  AOI21X1_65
timestamp 1522732896
transform 1 0 1880 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_177
timestamp 1522732896
transform -1 0 2008 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_29
timestamp 1522732896
transform 1 0 2008 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_367
timestamp 1522732896
transform 1 0 2040 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_114
timestamp 1522732896
transform 1 0 2104 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_108
timestamp 1522732896
transform -1 0 2360 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_370
timestamp 1522732896
transform -1 0 2424 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_124
timestamp 1522732896
transform 1 0 2424 0 -1 2610
box 0 0 32 200
use INVX4  INVX4_7
timestamp 1522732896
transform -1 0 2504 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_78
timestamp 1522732896
transform 1 0 2504 0 -1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_44
timestamp 1522732896
transform 1 0 2568 0 -1 2610
box 0 0 80 200
use INVX2  INVX2_24
timestamp 1522732896
transform 1 0 2648 0 -1 2610
box 0 0 32 200
use INVX2  INVX2_2
timestamp 1522732896
transform -1 0 2712 0 -1 2610
box 0 0 32 200
use AND2X2  AND2X2_39
timestamp 1522732896
transform 1 0 2712 0 -1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_33
timestamp 1522732896
transform 1 0 2776 0 -1 2610
box 0 0 80 200
use OAI22X1  OAI22X1_31
timestamp 1522732896
transform 1 0 2856 0 -1 2610
box 0 0 80 200
use AOI21X1  AOI21X1_66
timestamp 1522732896
transform 1 0 2936 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_59
timestamp 1522732896
transform -1 0 3064 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_173
timestamp 1522732896
transform 1 0 3064 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_1_0
timestamp 1522732896
transform 1 0 3128 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1522732896
transform 1 0 3144 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_2
timestamp 1522732896
transform 1 0 3160 0 -1 2610
box 0 0 16 200
use OAI22X1  OAI22X1_26
timestamp 1522732896
transform 1 0 3176 0 -1 2610
box 0 0 80 200
use AOI21X1  AOI21X1_58
timestamp 1522732896
transform -1 0 3320 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_62
timestamp 1522732896
transform 1 0 3320 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_90
timestamp 1522732896
transform 1 0 3384 0 -1 2610
box 0 0 192 200
use OAI22X1  OAI22X1_18
timestamp 1522732896
transform 1 0 3576 0 -1 2610
box 0 0 80 200
use INVX2  INVX2_42
timestamp 1522732896
transform -1 0 3688 0 -1 2610
box 0 0 32 200
use XNOR2X1  XNOR2X1_6
timestamp 1522732896
transform -1 0 3800 0 -1 2610
box 0 0 112 200
use NOR2X1  NOR2X1_227
timestamp 1522732896
transform 1 0 3800 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_148
timestamp 1522732896
transform 1 0 3848 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_224
timestamp 1522732896
transform -1 0 3944 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_164
timestamp 1522732896
transform 1 0 3944 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_225
timestamp 1522732896
transform 1 0 4008 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_270
timestamp 1522732896
transform 1 0 4056 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_269
timestamp 1522732896
transform 1 0 4120 0 -1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_4
timestamp 1522732896
transform -1 0 4280 0 -1 2610
box 0 0 96 200
use NAND2X1  NAND2X1_40
timestamp 1522732896
transform -1 0 4328 0 -1 2610
box 0 0 48 200
use AOI21X1  AOI21X1_38
timestamp 1522732896
transform 1 0 4328 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_64
timestamp 1522732896
transform -1 0 4456 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_273
timestamp 1522732896
transform 1 0 4456 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_43
timestamp 1522732896
transform -1 0 4584 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_33
timestamp 1522732896
transform -1 0 4616 0 -1 2610
box 0 0 32 200
use FILL  FILL_12_2_0
timestamp 1522732896
transform -1 0 4632 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1522732896
transform -1 0 4648 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_2
timestamp 1522732896
transform -1 0 4664 0 -1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_6
timestamp 1522732896
transform -1 0 4760 0 -1 2610
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_93
timestamp 1522732896
transform -1 0 4952 0 -1 2610
box 0 0 192 200
use AND2X2  AND2X2_40
timestamp 1522732896
transform -1 0 5016 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_57
timestamp 1522732896
transform -1 0 5208 0 -1 2610
box 0 0 192 200
use MUX2X1  MUX2X1_25
timestamp 1522732896
transform 1 0 5208 0 -1 2610
box 0 0 96 200
use INVX1  INVX1_148
timestamp 1522732896
transform -1 0 5336 0 -1 2610
box 0 0 32 200
use INVX1  INVX1_188
timestamp 1522732896
transform 1 0 5336 0 -1 2610
box 0 0 32 200
use AOI21X1  AOI21X1_127
timestamp 1522732896
transform 1 0 5368 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_58
timestamp 1522732896
transform 1 0 5432 0 -1 2610
box 0 0 80 200
use BUFX4  BUFX4_63
timestamp 1522732896
transform 1 0 5512 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_251
timestamp 1522732896
transform 1 0 5576 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_64
timestamp 1522732896
transform 1 0 5624 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_250
timestamp 1522732896
transform 1 0 5688 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_470
timestamp 1522732896
transform 1 0 5736 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_135
timestamp 1522732896
transform -1 0 5992 0 -1 2610
box 0 0 192 200
use INVX1  INVX1_189
timestamp 1522732896
transform 1 0 5992 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_472
timestamp 1522732896
transform 1 0 6024 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_137
timestamp 1522732896
transform -1 0 6280 0 -1 2610
box 0 0 192 200
use FILL  FILL_13_1
timestamp 1522732896
transform -1 0 6296 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_6
timestamp 1522732896
transform 1 0 8 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_122
timestamp 1522732896
transform 1 0 72 0 1 2210
box 0 0 192 200
use INVX2  INVX2_20
timestamp 1522732896
transform 1 0 264 0 1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_54
timestamp 1522732896
transform 1 0 296 0 1 2210
box 0 0 80 200
use NOR2X1  NOR2X1_223
timestamp 1522732896
transform -1 0 424 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_394
timestamp 1522732896
transform -1 0 488 0 1 2210
box 0 0 64 200
use INVX1  INVX1_162
timestamp 1522732896
transform -1 0 520 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_37
timestamp 1522732896
transform -1 0 584 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_37
timestamp 1522732896
transform -1 0 632 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_36
timestamp 1522732896
transform -1 0 680 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_38
timestamp 1522732896
transform 1 0 680 0 1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_33
timestamp 1522732896
transform 1 0 728 0 1 2210
box 0 0 64 200
use INVX1  INVX1_32
timestamp 1522732896
transform 1 0 792 0 1 2210
box 0 0 32 200
use NAND3X1  NAND3X1_42
timestamp 1522732896
transform 1 0 824 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_38
timestamp 1522732896
transform -1 0 936 0 1 2210
box 0 0 48 200
use OAI22X1  OAI22X1_5
timestamp 1522732896
transform -1 0 1016 0 1 2210
box 0 0 80 200
use INVX1  INVX1_8
timestamp 1522732896
transform 1 0 1016 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_123
timestamp 1522732896
transform 1 0 1048 0 1 2210
box 0 0 192 200
use INVX1  INVX1_1
timestamp 1522732896
transform 1 0 1240 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_41
timestamp 1522732896
transform -1 0 1336 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_4
timestamp 1522732896
transform -1 0 1400 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_38
timestamp 1522732896
transform 1 0 1400 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_41
timestamp 1522732896
transform -1 0 1528 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_12
timestamp 1522732896
transform 1 0 1528 0 1 2210
box 0 0 80 200
use FILL  FILL_11_0_0
timestamp 1522732896
transform -1 0 1624 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1522732896
transform -1 0 1640 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_2
timestamp 1522732896
transform -1 0 1656 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_42
timestamp 1522732896
transform -1 0 1720 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_35
timestamp 1522732896
transform -1 0 1784 0 1 2210
box 0 0 64 200
use INVX1  INVX1_31
timestamp 1522732896
transform 1 0 1784 0 1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_13
timestamp 1522732896
transform 1 0 1816 0 1 2210
box 0 0 48 200
use INVX1  INVX1_156
timestamp 1522732896
transform 1 0 1864 0 1 2210
box 0 0 32 200
use NAND3X1  NAND3X1_149
timestamp 1522732896
transform 1 0 1896 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_109
timestamp 1522732896
transform -1 0 2152 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_372
timestamp 1522732896
transform 1 0 2152 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_346
timestamp 1522732896
transform -1 0 2280 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_194
timestamp 1522732896
transform 1 0 2280 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_88
timestamp 1522732896
transform 1 0 2344 0 1 2210
box 0 0 192 200
use AOI21X1  AOI21X1_69
timestamp 1522732896
transform 1 0 2536 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_186
timestamp 1522732896
transform -1 0 2664 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_68
timestamp 1522732896
transform -1 0 2728 0 1 2210
box 0 0 64 200
use OAI22X1  OAI22X1_27
timestamp 1522732896
transform 1 0 2728 0 1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_168
timestamp 1522732896
transform -1 0 2872 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_147
timestamp 1522732896
transform -1 0 2920 0 1 2210
box 0 0 48 200
use INVX1  INVX1_114
timestamp 1522732896
transform 1 0 2920 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_181
timestamp 1522732896
transform -1 0 3016 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_76
timestamp 1522732896
transform -1 0 3208 0 1 2210
box 0 0 192 200
use FILL  FILL_11_1_0
timestamp 1522732896
transform -1 0 3224 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1522732896
transform -1 0 3240 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_2
timestamp 1522732896
transform -1 0 3256 0 1 2210
box 0 0 16 200
use BUFX2  BUFX2_10
timestamp 1522732896
transform -1 0 3304 0 1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_87
timestamp 1522732896
transform -1 0 3368 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_42
timestamp 1522732896
transform -1 0 3448 0 1 2210
box 0 0 80 200
use INVX1  INVX1_151
timestamp 1522732896
transform -1 0 3480 0 1 2210
box 0 0 32 200
use AND2X2  AND2X2_44
timestamp 1522732896
transform -1 0 3544 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_297
timestamp 1522732896
transform 1 0 3544 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_86
timestamp 1522732896
transform 1 0 3608 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_84
timestamp 1522732896
transform 1 0 3672 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_179
timestamp 1522732896
transform 1 0 3736 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_282
timestamp 1522732896
transform -1 0 3848 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_26
timestamp 1522732896
transform -1 0 3944 0 1 2210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_87
timestamp 1522732896
transform 1 0 3944 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_281
timestamp 1522732896
transform 1 0 4136 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_21
timestamp 1522732896
transform -1 0 4264 0 1 2210
box 0 0 64 200
use INVX2  INVX2_33
timestamp 1522732896
transform -1 0 4296 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_268
timestamp 1522732896
transform 1 0 4296 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_267
timestamp 1522732896
transform 1 0 4360 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_133
timestamp 1522732896
transform -1 0 4488 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_134
timestamp 1522732896
transform 1 0 4488 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_77
timestamp 1522732896
transform -1 0 4744 0 1 2210
box 0 0 192 200
use FILL  FILL_11_2_0
timestamp 1522732896
transform 1 0 4744 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1522732896
transform 1 0 4760 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_2
timestamp 1522732896
transform 1 0 4776 0 1 2210
box 0 0 16 200
use INVX1  INVX1_116
timestamp 1522732896
transform 1 0 4792 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_56
timestamp 1522732896
transform -1 0 5016 0 1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_85
timestamp 1522732896
transform 1 0 5016 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_46
timestamp 1522732896
transform 1 0 5208 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_84
timestamp 1522732896
transform -1 0 5448 0 1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_136
timestamp 1522732896
transform -1 0 5640 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_471
timestamp 1522732896
transform -1 0 5704 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_212
timestamp 1522732896
transform 1 0 5704 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_458
timestamp 1522732896
transform -1 0 5816 0 1 2210
box 0 0 64 200
use XNOR2X1  XNOR2X1_9
timestamp 1522732896
transform 1 0 5816 0 1 2210
box 0 0 112 200
use OAI21X1  OAI21X1_473
timestamp 1522732896
transform 1 0 5928 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_253
timestamp 1522732896
transform -1 0 6040 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_138
timestamp 1522732896
transform -1 0 6232 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_459
timestamp 1522732896
transform 1 0 6232 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_116
timestamp 1522732896
transform -1 0 200 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_384
timestamp 1522732896
transform -1 0 264 0 -1 2210
box 0 0 64 200
use INVX2  INVX2_7
timestamp 1522732896
transform 1 0 264 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_382
timestamp 1522732896
transform 1 0 296 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_5
timestamp 1522732896
transform 1 0 360 0 -1 2210
box 0 0 80 200
use NAND3X1  NAND3X1_15
timestamp 1522732896
transform 1 0 440 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_124
timestamp 1522732896
transform 1 0 504 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_40
timestamp 1522732896
transform 1 0 696 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_37
timestamp 1522732896
transform -1 0 808 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_7
timestamp 1522732896
transform 1 0 808 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_26
timestamp 1522732896
transform -1 0 936 0 -1 2210
box 0 0 80 200
use NAND3X1  NAND3X1_13
timestamp 1522732896
transform -1 0 1000 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_14
timestamp 1522732896
transform 1 0 1000 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_29
timestamp 1522732896
transform -1 0 1144 0 -1 2210
box 0 0 80 200
use BUFX2  BUFX2_12
timestamp 1522732896
transform -1 0 1192 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_12
timestamp 1522732896
transform -1 0 1256 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_20
timestamp 1522732896
transform 1 0 1256 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_12
timestamp 1522732896
transform -1 0 1352 0 -1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_12
timestamp 1522732896
transform 1 0 1352 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_18
timestamp 1522732896
transform 1 0 1416 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_16
timestamp 1522732896
transform -1 0 1528 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_10
timestamp 1522732896
transform -1 0 1592 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_0_0
timestamp 1522732896
transform -1 0 1608 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1522732896
transform -1 0 1624 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_2
timestamp 1522732896
transform -1 0 1640 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_13
timestamp 1522732896
transform -1 0 1704 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_21
timestamp 1522732896
transform -1 0 1752 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_28
timestamp 1522732896
transform -1 0 1832 0 -1 2210
box 0 0 80 200
use INVX2  INVX2_8
timestamp 1522732896
transform -1 0 1864 0 -1 2210
box 0 0 32 200
use INVX2  INVX2_38
timestamp 1522732896
transform -1 0 1896 0 -1 2210
box 0 0 32 200
use INVX8  INVX8_4
timestamp 1522732896
transform 1 0 1896 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_4
timestamp 1522732896
transform -1 0 2040 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_76
timestamp 1522732896
transform 1 0 2040 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_15
timestamp 1522732896
transform -1 0 2168 0 -1 2210
box 0 0 64 200
use INVX2  INVX2_34
timestamp 1522732896
transform -1 0 2200 0 -1 2210
box 0 0 32 200
use INVX2  INVX2_36
timestamp 1522732896
transform -1 0 2232 0 -1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_195
timestamp 1522732896
transform 1 0 2232 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_190
timestamp 1522732896
transform 1 0 2280 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_36
timestamp 1522732896
transform 1 0 2344 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_139
timestamp 1522732896
transform -1 0 2472 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_17
timestamp 1522732896
transform 1 0 2472 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_150
timestamp 1522732896
transform -1 0 2584 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_185
timestamp 1522732896
transform -1 0 2648 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_184
timestamp 1522732896
transform -1 0 2712 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_61
timestamp 1522732896
transform 1 0 2712 0 -1 2210
box 0 0 64 200
use INVX2  INVX2_37
timestamp 1522732896
transform -1 0 2808 0 -1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_28
timestamp 1522732896
transform 1 0 2808 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_169
timestamp 1522732896
transform -1 0 2952 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_179
timestamp 1522732896
transform -1 0 3016 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_3
timestamp 1522732896
transform 1 0 3016 0 -1 2210
box 0 0 96 200
use FILL  FILL_10_1_0
timestamp 1522732896
transform 1 0 3112 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1522732896
transform 1 0 3128 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_2
timestamp 1522732896
transform 1 0 3144 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_298
timestamp 1522732896
transform 1 0 3160 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_115
timestamp 1522732896
transform -1 0 3256 0 -1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_89
timestamp 1522732896
transform -1 0 3448 0 -1 2210
box 0 0 192 200
use AOI22X1  AOI22X1_41
timestamp 1522732896
transform -1 0 3528 0 -1 2210
box 0 0 80 200
use INVX1  INVX1_46
timestamp 1522732896
transform 1 0 3528 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_296
timestamp 1522732896
transform 1 0 3560 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_292
timestamp 1522732896
transform 1 0 3624 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_293
timestamp 1522732896
transform -1 0 3752 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_83
timestamp 1522732896
transform -1 0 3816 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_189
timestamp 1522732896
transform -1 0 3864 0 -1 2210
box 0 0 48 200
use OAI22X1  OAI22X1_42
timestamp 1522732896
transform 1 0 3864 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_303
timestamp 1522732896
transform 1 0 3944 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_91
timestamp 1522732896
transform 1 0 4008 0 -1 2210
box 0 0 192 200
use AOI21X1  AOI21X1_88
timestamp 1522732896
transform -1 0 4264 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_125
timestamp 1522732896
transform 1 0 4264 0 -1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_45
timestamp 1522732896
transform 1 0 4296 0 -1 2210
box 0 0 48 200
use MUX2X1  MUX2X1_5
timestamp 1522732896
transform -1 0 4440 0 -1 2210
box 0 0 96 200
use OAI21X1  OAI21X1_84
timestamp 1522732896
transform 1 0 4440 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_40
timestamp 1522732896
transform -1 0 4568 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_43
timestamp 1522732896
transform -1 0 4600 0 -1 2210
box 0 0 32 200
use INVX4  INVX4_2
timestamp 1522732896
transform 1 0 4600 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_2_0
timestamp 1522732896
transform 1 0 4648 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1522732896
transform 1 0 4664 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_2
timestamp 1522732896
transform 1 0 4680 0 -1 2210
box 0 0 16 200
use INVX1  INVX1_60
timestamp 1522732896
transform 1 0 4696 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_280
timestamp 1522732896
transform 1 0 4728 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_188
timestamp 1522732896
transform 1 0 4792 0 -1 2210
box 0 0 48 200
use INVX2  INVX2_43
timestamp 1522732896
transform -1 0 4872 0 -1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_39
timestamp 1522732896
transform 1 0 4872 0 -1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_163
timestamp 1522732896
transform -1 0 5000 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_149
timestamp 1522732896
transform 1 0 5000 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_45
timestamp 1522732896
transform 1 0 5048 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_44
timestamp 1522732896
transform 1 0 5112 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_150
timestamp 1522732896
transform -1 0 5192 0 -1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_42
timestamp 1522732896
transform -1 0 5384 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_43
timestamp 1522732896
transform -1 0 5576 0 -1 2210
box 0 0 192 200
use INVX2  INVX2_31
timestamp 1522732896
transform -1 0 5608 0 -1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_126
timestamp 1522732896
transform -1 0 5800 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_23
timestamp 1522732896
transform 1 0 5800 0 -1 2210
box 0 0 64 200
use XNOR2X1  XNOR2X1_10
timestamp 1522732896
transform -1 0 5976 0 -1 2210
box 0 0 112 200
use XOR2X1  XOR2X1_3
timestamp 1522732896
transform -1 0 6088 0 -1 2210
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_127
timestamp 1522732896
transform -1 0 6280 0 -1 2210
box 0 0 192 200
use FILL  FILL_11_1
timestamp 1522732896
transform -1 0 6296 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_117
timestamp 1522732896
transform -1 0 200 0 1 1810
box 0 0 192 200
use AOI21X1  AOI21X1_118
timestamp 1522732896
transform 1 0 200 0 1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_50
timestamp 1522732896
transform -1 0 344 0 1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_385
timestamp 1522732896
transform 1 0 344 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_12
timestamp 1522732896
transform 1 0 408 0 1 1810
box 0 0 64 200
use INVX2  INVX2_6
timestamp 1522732896
transform 1 0 472 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_206
timestamp 1522732896
transform 1 0 504 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_17
timestamp 1522732896
transform -1 0 616 0 1 1810
box 0 0 64 200
use INVX1  INVX1_157
timestamp 1522732896
transform 1 0 616 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_375
timestamp 1522732896
transform -1 0 712 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_373
timestamp 1522732896
transform -1 0 776 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_68
timestamp 1522732896
transform 1 0 776 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_183
timestamp 1522732896
transform -1 0 1032 0 1 1810
box 0 0 64 200
use INVX1  INVX1_117
timestamp 1522732896
transform -1 0 1064 0 1 1810
box 0 0 32 200
use AOI21X1  AOI21X1_9
timestamp 1522732896
transform -1 0 1128 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_374
timestamp 1522732896
transform 1 0 1128 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1522732896
transform -1 0 1256 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1522732896
transform 1 0 1256 0 1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_1
timestamp 1522732896
transform 1 0 1320 0 1 1810
box 0 0 80 200
use AOI21X1  AOI21X1_13
timestamp 1522732896
transform -1 0 1464 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_15
timestamp 1522732896
transform 1 0 1464 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_27
timestamp 1522732896
transform 1 0 1528 0 1 1810
box 0 0 64 200
use FILL  FILL_9_0_0
timestamp 1522732896
transform 1 0 1592 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1522732896
transform 1 0 1608 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_2
timestamp 1522732896
transform 1 0 1624 0 1 1810
box 0 0 16 200
use INVX4  INVX4_1
timestamp 1522732896
transform 1 0 1640 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_213
timestamp 1522732896
transform -1 0 1736 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_81
timestamp 1522732896
transform 1 0 1736 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_28
timestamp 1522732896
transform 1 0 1800 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_202
timestamp 1522732896
transform -1 0 1912 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_204
timestamp 1522732896
transform 1 0 1912 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_153
timestamp 1522732896
transform 1 0 1960 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_161
timestamp 1522732896
transform 1 0 2024 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_138
timestamp 1522732896
transform 1 0 2088 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_193
timestamp 1522732896
transform 1 0 2152 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_144
timestamp 1522732896
transform 1 0 2200 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_194
timestamp 1522732896
transform -1 0 2296 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_148
timestamp 1522732896
transform -1 0 2360 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_135
timestamp 1522732896
transform 1 0 2360 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_72
timestamp 1522732896
transform -1 0 2472 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_71
timestamp 1522732896
transform -1 0 2536 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_79
timestamp 1522732896
transform 1 0 2536 0 1 1810
box 0 0 64 200
use INVX1  INVX1_65
timestamp 1522732896
transform 1 0 2600 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_131
timestamp 1522732896
transform -1 0 2680 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_93
timestamp 1522732896
transform 1 0 2680 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_136
timestamp 1522732896
transform 1 0 2744 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_92
timestamp 1522732896
transform 1 0 2792 0 1 1810
box 0 0 64 200
use INVX4  INVX4_4
timestamp 1522732896
transform 1 0 2856 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_187
timestamp 1522732896
transform 1 0 2904 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_145
timestamp 1522732896
transform 1 0 2952 0 1 1810
box 0 0 48 200
use INVX2  INVX2_40
timestamp 1522732896
transform 1 0 3000 0 1 1810
box 0 0 32 200
use MUX2X1  MUX2X1_10
timestamp 1522732896
transform 1 0 3032 0 1 1810
box 0 0 96 200
use FILL  FILL_9_1_0
timestamp 1522732896
transform 1 0 3128 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1522732896
transform 1 0 3144 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_2
timestamp 1522732896
transform 1 0 3160 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_278
timestamp 1522732896
transform 1 0 3176 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_178
timestamp 1522732896
transform 1 0 3240 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_190
timestamp 1522732896
transform 1 0 3288 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_295
timestamp 1522732896
transform 1 0 3336 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_186
timestamp 1522732896
transform -1 0 3448 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_85
timestamp 1522732896
transform -1 0 3512 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_294
timestamp 1522732896
transform -1 0 3576 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_99
timestamp 1522732896
transform -1 0 3624 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_17
timestamp 1522732896
transform -1 0 3688 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_146
timestamp 1522732896
transform -1 0 3752 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_291
timestamp 1522732896
transform -1 0 3816 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_302
timestamp 1522732896
transform 1 0 3816 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_189
timestamp 1522732896
transform -1 0 3928 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_191
timestamp 1522732896
transform 1 0 3928 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_70
timestamp 1522732896
transform 1 0 3976 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_300
timestamp 1522732896
transform 1 0 4040 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_301
timestamp 1522732896
transform -1 0 4168 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_272
timestamp 1522732896
transform 1 0 4168 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_271
timestamp 1522732896
transform 1 0 4232 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_42
timestamp 1522732896
transform -1 0 4344 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_79
timestamp 1522732896
transform -1 0 4536 0 1 1810
box 0 0 192 200
use AOI21X1  AOI21X1_82
timestamp 1522732896
transform 1 0 4536 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_147
timestamp 1522732896
transform 1 0 4600 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1522732896
transform 1 0 4664 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1522732896
transform 1 0 4680 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_2
timestamp 1522732896
transform 1 0 4696 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_81
timestamp 1522732896
transform 1 0 4712 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_185
timestamp 1522732896
transform -1 0 4824 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_277
timestamp 1522732896
transform -1 0 4888 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_231
timestamp 1522732896
transform 1 0 4888 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_136
timestamp 1522732896
transform -1 0 5016 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_276
timestamp 1522732896
transform 1 0 5016 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_275
timestamp 1522732896
transform -1 0 5144 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_46
timestamp 1522732896
transform 1 0 5144 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_207
timestamp 1522732896
transform -1 0 5272 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_209
timestamp 1522732896
transform 1 0 5272 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_208
timestamp 1522732896
transform -1 0 5400 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_210
timestamp 1522732896
transform -1 0 5464 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_44
timestamp 1522732896
transform -1 0 5656 0 1 1810
box 0 0 192 200
use BUFX4  BUFX4_25
timestamp 1522732896
transform -1 0 5720 0 1 1810
box 0 0 64 200
use INVX1  INVX1_119
timestamp 1522732896
transform -1 0 5752 0 1 1810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_45
timestamp 1522732896
transform 1 0 5752 0 1 1810
box 0 0 192 200
use INVX1  INVX1_105
timestamp 1522732896
transform 1 0 5944 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_146
timestamp 1522732896
transform -1 0 6024 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_163
timestamp 1522732896
transform -1 0 6088 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_162
timestamp 1522732896
transform 1 0 6088 0 1 1810
box 0 0 64 200
use INVX1  INVX1_104
timestamp 1522732896
transform -1 0 6184 0 1 1810
box 0 0 32 200
use INVX1  INVX1_195
timestamp 1522732896
transform -1 0 6216 0 1 1810
box 0 0 32 200
use OR2X2  OR2X2_41
timestamp 1522732896
transform -1 0 6280 0 1 1810
box 0 0 64 200
use FILL  FILL_10_1
timestamp 1522732896
transform 1 0 6280 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_117
timestamp 1522732896
transform 1 0 8 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_383
timestamp 1522732896
transform -1 0 136 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_161
timestamp 1522732896
transform -1 0 200 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_209
timestamp 1522732896
transform -1 0 248 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_110
timestamp 1522732896
transform 1 0 248 0 -1 1810
box 0 0 192 200
use INVX2  INVX2_9
timestamp 1522732896
transform 1 0 440 0 -1 1810
box 0 0 32 200
use OAI22X1  OAI22X1_45
timestamp 1522732896
transform 1 0 472 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_215
timestamp 1522732896
transform 1 0 552 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_6
timestamp 1522732896
transform -1 0 680 0 -1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_205
timestamp 1522732896
transform -1 0 728 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_24
timestamp 1522732896
transform -1 0 776 0 -1 1810
box 0 0 48 200
use NOR3X1  NOR3X1_3
timestamp 1522732896
transform 1 0 776 0 -1 1810
box 0 0 128 200
use BUFX4  BUFX4_82
timestamp 1522732896
transform 1 0 904 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_70
timestamp 1522732896
transform -1 0 1032 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_4
timestamp 1522732896
transform 1 0 1032 0 -1 1810
box 0 0 80 200
use BUFX4  BUFX4_80
timestamp 1522732896
transform -1 0 1176 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_31
timestamp 1522732896
transform 1 0 1176 0 -1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_2
timestamp 1522732896
transform -1 0 1320 0 -1 1810
box 0 0 80 200
use BUFX4  BUFX4_72
timestamp 1522732896
transform 1 0 1320 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_134
timestamp 1522732896
transform 1 0 1384 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_201
timestamp 1522732896
transform -1 0 1496 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_152
timestamp 1522732896
transform 1 0 1496 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1522732896
transform -1 0 1576 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1522732896
transform -1 0 1592 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_2
timestamp 1522732896
transform -1 0 1608 0 -1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_92
timestamp 1522732896
transform -1 0 1672 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_14
timestamp 1522732896
transform 1 0 1672 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_203
timestamp 1522732896
transform 1 0 1736 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_155
timestamp 1522732896
transform 1 0 1784 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_132
timestamp 1522732896
transform 1 0 1848 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_196
timestamp 1522732896
transform 1 0 1896 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_122
timestamp 1522732896
transform 1 0 1944 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_208
timestamp 1522732896
transform -1 0 2040 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_43
timestamp 1522732896
transform 1 0 2040 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_188
timestamp 1522732896
transform 1 0 2104 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_151
timestamp 1522732896
transform -1 0 2216 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_195
timestamp 1522732896
transform -1 0 2264 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_314
timestamp 1522732896
transform 1 0 2264 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_205
timestamp 1522732896
transform -1 0 2376 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_123
timestamp 1522732896
transform 1 0 2376 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_134
timestamp 1522732896
transform -1 0 2472 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_141
timestamp 1522732896
transform -1 0 2520 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_142
timestamp 1522732896
transform 1 0 2520 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_102
timestamp 1522732896
transform -1 0 2632 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_143
timestamp 1522732896
transform -1 0 2680 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_230
timestamp 1522732896
transform 1 0 2680 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_130
timestamp 1522732896
transform -1 0 2792 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_91
timestamp 1522732896
transform -1 0 2856 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_64
timestamp 1522732896
transform -1 0 2888 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_121
timestamp 1522732896
transform -1 0 2936 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_142
timestamp 1522732896
transform 1 0 2936 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_75
timestamp 1522732896
transform -1 0 3176 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_1_0
timestamp 1522732896
transform 1 0 3176 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1522732896
transform 1 0 3192 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_2
timestamp 1522732896
transform 1 0 3208 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_266
timestamp 1522732896
transform 1 0 3224 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_40
timestamp 1522732896
transform -1 0 3368 0 -1 1810
box 0 0 80 200
use INVX1  INVX1_139
timestamp 1522732896
transform 1 0 3368 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_108
timestamp 1522732896
transform 1 0 3400 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_164
timestamp 1522732896
transform 1 0 3432 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_60
timestamp 1522732896
transform -1 0 3560 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_91
timestamp 1522732896
transform 1 0 3560 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_92
timestamp 1522732896
transform 1 0 3624 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_100
timestamp 1522732896
transform 1 0 3688 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_191
timestamp 1522732896
transform 1 0 3736 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_42
timestamp 1522732896
transform -1 0 3848 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_279
timestamp 1522732896
transform -1 0 3912 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_86
timestamp 1522732896
transform 1 0 3912 0 -1 1810
box 0 0 192 200
use INVX2  INVX2_28
timestamp 1522732896
transform 1 0 4104 0 -1 1810
box 0 0 32 200
use BUFX4  BUFX4_36
timestamp 1522732896
transform -1 0 4200 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_44
timestamp 1522732896
transform 1 0 4200 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_24
timestamp 1522732896
transform 1 0 4264 0 -1 1810
box 0 0 96 200
use INVX1  INVX1_147
timestamp 1522732896
transform -1 0 4392 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_85
timestamp 1522732896
transform 1 0 4392 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_83
timestamp 1522732896
transform 1 0 4456 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_2_0
timestamp 1522732896
transform 1 0 4648 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1522732896
transform 1 0 4664 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_2
timestamp 1522732896
transform 1 0 4680 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_299
timestamp 1522732896
transform 1 0 4696 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_190
timestamp 1522732896
transform 1 0 4760 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_130
timestamp 1522732896
transform -1 0 4872 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_164
timestamp 1522732896
transform -1 0 4920 0 -1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_51
timestamp 1522732896
transform -1 0 4984 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_50
timestamp 1522732896
transform -1 0 5048 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_61
timestamp 1522732896
transform -1 0 5080 0 -1 1810
box 0 0 32 200
use BUFX4  BUFX4_44
timestamp 1522732896
transform 1 0 5080 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_202
timestamp 1522732896
transform 1 0 5144 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_204
timestamp 1522732896
transform -1 0 5272 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_40
timestamp 1522732896
transform -1 0 5464 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_211
timestamp 1522732896
transform 1 0 5464 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_212
timestamp 1522732896
transform -1 0 5592 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_156
timestamp 1522732896
transform -1 0 5640 0 -1 1810
box 0 0 48 200
use OAI22X1  OAI22X1_36
timestamp 1522732896
transform -1 0 5720 0 -1 1810
box 0 0 80 200
use INVX1  INVX1_132
timestamp 1522732896
transform 1 0 5720 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_206
timestamp 1522732896
transform 1 0 5752 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_205
timestamp 1522732896
transform 1 0 5816 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_47
timestamp 1522732896
transform -1 0 6072 0 -1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_41
timestamp 1522732896
transform -1 0 6264 0 -1 1810
box 0 0 192 200
use FILL  FILL_9_1
timestamp 1522732896
transform -1 0 6280 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_2
timestamp 1522732896
transform -1 0 6296 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_27
timestamp 1522732896
transform -1 0 72 0 1 1410
box 0 0 64 200
use INVX1  INVX1_23
timestamp 1522732896
transform -1 0 104 0 1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_70
timestamp 1522732896
transform -1 0 296 0 1 1410
box 0 0 192 200
use INVX4  INVX4_6
timestamp 1522732896
transform 1 0 296 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_22
timestamp 1522732896
transform -1 0 408 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_137
timestamp 1522732896
transform 1 0 408 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_83
timestamp 1522732896
transform -1 0 536 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_10
timestamp 1522732896
transform -1 0 584 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_4
timestamp 1522732896
transform 1 0 584 0 1 1410
box 0 0 64 200
use INVX1  INVX1_15
timestamp 1522732896
transform 1 0 648 0 1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_11
timestamp 1522732896
transform -1 0 728 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_16
timestamp 1522732896
transform 1 0 728 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_196
timestamp 1522732896
transform -1 0 840 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_152
timestamp 1522732896
transform -1 0 904 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1522732896
transform 1 0 904 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_66
timestamp 1522732896
transform 1 0 952 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_151
timestamp 1522732896
transform -1 0 1064 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_27
timestamp 1522732896
transform 1 0 1064 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_193
timestamp 1522732896
transform 1 0 1128 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_150
timestamp 1522732896
transform -1 0 1240 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_158
timestamp 1522732896
transform 1 0 1240 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_45
timestamp 1522732896
transform -1 0 1368 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_309
timestamp 1522732896
transform 1 0 1368 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_212
timestamp 1522732896
transform 1 0 1432 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_210
timestamp 1522732896
transform -1 0 1528 0 1 1410
box 0 0 48 200
use INVX1  INVX1_154
timestamp 1522732896
transform -1 0 1560 0 1 1410
box 0 0 32 200
use FILL  FILL_7_0_0
timestamp 1522732896
transform -1 0 1576 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1522732896
transform -1 0 1592 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_2
timestamp 1522732896
transform -1 0 1608 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_310
timestamp 1522732896
transform -1 0 1672 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_129
timestamp 1522732896
transform 1 0 1672 0 1 1410
box 0 0 64 200
use INVX1  INVX1_62
timestamp 1522732896
transform 1 0 1736 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_306
timestamp 1522732896
transform -1 0 1832 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_197
timestamp 1522732896
transform -1 0 1880 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_74
timestamp 1522732896
transform 1 0 1880 0 1 1410
box 0 0 48 200
use INVX1  INVX1_39
timestamp 1522732896
transform -1 0 1960 0 1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_154
timestamp 1522732896
transform -1 0 2024 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_14
timestamp 1522732896
transform -1 0 2152 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_187
timestamp 1522732896
transform 1 0 2152 0 1 1410
box 0 0 64 200
use INVX1  INVX1_153
timestamp 1522732896
transform 1 0 2216 0 1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_92
timestamp 1522732896
transform -1 0 2296 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_145
timestamp 1522732896
transform -1 0 2360 0 1 1410
box 0 0 64 200
use INVX1  INVX1_118
timestamp 1522732896
transform 1 0 2360 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_1
timestamp 1522732896
transform 1 0 2392 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_101
timestamp 1522732896
transform -1 0 2520 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_139
timestamp 1522732896
transform 1 0 2520 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_95
timestamp 1522732896
transform -1 0 2632 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_12
timestamp 1522732896
transform 1 0 2632 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_165
timestamp 1522732896
transform -1 0 2824 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_140
timestamp 1522732896
transform 1 0 2824 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_148
timestamp 1522732896
transform 1 0 2872 0 1 1410
box 0 0 64 200
use INVX1  INVX1_112
timestamp 1522732896
transform 1 0 2936 0 1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_96
timestamp 1522732896
transform -1 0 3032 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_125
timestamp 1522732896
transform -1 0 3080 0 1 1410
box 0 0 48 200
use FILL  FILL_7_1_0
timestamp 1522732896
transform 1 0 3080 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1522732896
transform 1 0 3096 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_2
timestamp 1522732896
transform 1 0 3112 0 1 1410
box 0 0 16 200
use MUX2X1  MUX2X1_2
timestamp 1522732896
transform 1 0 3128 0 1 1410
box 0 0 96 200
use OAI21X1  OAI21X1_304
timestamp 1522732896
transform -1 0 3288 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_92
timestamp 1522732896
transform 1 0 3288 0 1 1410
box 0 0 192 200
use INVX1  INVX1_107
timestamp 1522732896
transform 1 0 3480 0 1 1410
box 0 0 32 200
use XNOR2X1  XNOR2X1_1
timestamp 1522732896
transform 1 0 3512 0 1 1410
box 0 0 112 200
use MUX2X1  MUX2X1_9
timestamp 1522732896
transform -1 0 3720 0 1 1410
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_37
timestamp 1522732896
transform -1 0 3912 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_153
timestamp 1522732896
transform 1 0 3912 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_201
timestamp 1522732896
transform -1 0 4024 0 1 1410
box 0 0 64 200
use INVX2  INVX2_39
timestamp 1522732896
transform 1 0 4024 0 1 1410
box 0 0 32 200
use BUFX4  BUFX4_16
timestamp 1522732896
transform 1 0 4056 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_146
timestamp 1522732896
transform -1 0 4184 0 1 1410
box 0 0 64 200
use INVX1  INVX1_69
timestamp 1522732896
transform 1 0 4184 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_147
timestamp 1522732896
transform -1 0 4280 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_73
timestamp 1522732896
transform 1 0 4280 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_84
timestamp 1522732896
transform 1 0 4344 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_35
timestamp 1522732896
transform -1 0 4584 0 1 1410
box 0 0 192 200
use INVX2  INVX2_32
timestamp 1522732896
transform 1 0 4584 0 1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_90
timestamp 1522732896
transform -1 0 4680 0 1 1410
box 0 0 64 200
use FILL  FILL_7_2_0
timestamp 1522732896
transform 1 0 4680 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1522732896
transform 1 0 4696 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_2
timestamp 1522732896
transform 1 0 4712 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_151
timestamp 1522732896
transform 1 0 4728 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_199
timestamp 1522732896
transform -1 0 4840 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_129
timestamp 1522732896
transform 1 0 4840 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_71
timestamp 1522732896
transform -1 0 4952 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_13
timestamp 1522732896
transform -1 0 5016 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_45
timestamp 1522732896
transform 1 0 5016 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_52
timestamp 1522732896
transform -1 0 5272 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_225
timestamp 1522732896
transform -1 0 5336 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_226
timestamp 1522732896
transform -1 0 5400 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_18
timestamp 1522732896
transform 1 0 5400 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_58
timestamp 1522732896
transform -1 0 5656 0 1 1410
box 0 0 192 200
use BUFX4  BUFX4_41
timestamp 1522732896
transform 1 0 5656 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_243
timestamp 1522732896
transform 1 0 5720 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_223
timestamp 1522732896
transform 1 0 5784 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_228
timestamp 1522732896
transform 1 0 5848 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_217
timestamp 1522732896
transform 1 0 5912 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_224
timestamp 1522732896
transform -1 0 6040 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_218
timestamp 1522732896
transform -1 0 6104 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_50
timestamp 1522732896
transform -1 0 6296 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_30
timestamp 1522732896
transform -1 0 56 0 -1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_2
timestamp 1522732896
transform -1 0 184 0 -1 1410
box 0 0 128 200
use NOR2X1  NOR2X1_133
timestamp 1522732896
transform 1 0 184 0 -1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_1
timestamp 1522732896
transform -1 0 360 0 -1 1410
box 0 0 128 200
use NOR2X1  NOR2X1_14
timestamp 1522732896
transform -1 0 408 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_17
timestamp 1522732896
transform -1 0 456 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_85
timestamp 1522732896
transform -1 0 520 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1522732896
transform 1 0 520 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_7
timestamp 1522732896
transform 1 0 584 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_2
timestamp 1522732896
transform 1 0 648 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_16
timestamp 1522732896
transform 1 0 712 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_17
timestamp 1522732896
transform 1 0 744 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_22
timestamp 1522732896
transform -1 0 856 0 -1 1410
box 0 0 48 200
use INVX8  INVX8_2
timestamp 1522732896
transform -1 0 936 0 -1 1410
box 0 0 80 200
use OAI22X1  OAI22X1_7
timestamp 1522732896
transform 1 0 936 0 -1 1410
box 0 0 80 200
use INVX1  INVX1_48
timestamp 1522732896
transform 1 0 1016 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_151
timestamp 1522732896
transform -1 0 1112 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_102
timestamp 1522732896
transform -1 0 1160 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_313
timestamp 1522732896
transform 1 0 1160 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_10
timestamp 1522732896
transform 1 0 1224 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_198
timestamp 1522732896
transform 1 0 1288 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_209
timestamp 1522732896
transform -1 0 1384 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_79
timestamp 1522732896
transform 1 0 1384 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_124
timestamp 1522732896
transform 1 0 1432 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_189
timestamp 1522732896
transform -1 0 1544 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_133
timestamp 1522732896
transform 1 0 1544 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_0_0
timestamp 1522732896
transform -1 0 1624 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1522732896
transform -1 0 1640 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_2
timestamp 1522732896
transform -1 0 1656 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_307
timestamp 1522732896
transform -1 0 1720 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_305
timestamp 1522732896
transform -1 0 1784 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_87
timestamp 1522732896
transform -1 0 1848 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_22
timestamp 1522732896
transform 1 0 1848 0 -1 1410
box 0 0 64 200
use OAI22X1  OAI22X1_20
timestamp 1522732896
transform 1 0 1912 0 -1 1410
box 0 0 80 200
use BUFX4  BUFX4_48
timestamp 1522732896
transform -1 0 2056 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_49
timestamp 1522732896
transform 1 0 2056 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_63
timestamp 1522732896
transform -1 0 2152 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_144
timestamp 1522732896
transform 1 0 2152 0 -1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_13
timestamp 1522732896
transform -1 0 2344 0 -1 1410
box 0 0 128 200
use BUFX4  BUFX4_86
timestamp 1522732896
transform 1 0 2344 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_135
timestamp 1522732896
transform 1 0 2408 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_11
timestamp 1522732896
transform 1 0 2472 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_143
timestamp 1522732896
transform -1 0 2600 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_51
timestamp 1522732896
transform -1 0 2648 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_46
timestamp 1522732896
transform 1 0 2648 0 -1 1410
box 0 0 64 200
use OAI22X1  OAI22X1_19
timestamp 1522732896
transform 1 0 2712 0 -1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_140
timestamp 1522732896
transform 1 0 2792 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_131
timestamp 1522732896
transform 1 0 2856 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_132
timestamp 1522732896
transform 1 0 2920 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_149
timestamp 1522732896
transform 1 0 2984 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_96
timestamp 1522732896
transform -1 0 3096 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_111
timestamp 1522732896
transform 1 0 3096 0 -1 1410
box 0 0 32 200
use FILL  FILL_6_1_0
timestamp 1522732896
transform 1 0 3128 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1522732896
transform 1 0 3144 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_2
timestamp 1522732896
transform 1 0 3160 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_9
timestamp 1522732896
transform 1 0 3176 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_192
timestamp 1522732896
transform -1 0 3288 0 -1 1410
box 0 0 48 200
use XOR2X1  XOR2X1_1
timestamp 1522732896
transform 1 0 3288 0 -1 1410
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_65
timestamp 1522732896
transform -1 0 3592 0 -1 1410
box 0 0 192 200
use NOR2X1  NOR2X1_152
timestamp 1522732896
transform -1 0 3640 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_144
timestamp 1522732896
transform 1 0 3640 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_259
timestamp 1522732896
transform 1 0 3672 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_63
timestamp 1522732896
transform 1 0 3736 0 -1 1410
box 0 0 192 200
use INVX1  INVX1_141
timestamp 1522732896
transform 1 0 3928 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_251
timestamp 1522732896
transform 1 0 3960 0 -1 1410
box 0 0 64 200
use OAI22X1  OAI22X1_35
timestamp 1522732896
transform 1 0 4024 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_39
timestamp 1522732896
transform -1 0 4296 0 -1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_176
timestamp 1522732896
transform 1 0 4296 0 -1 1410
box 0 0 48 200
use OAI22X1  OAI22X1_34
timestamp 1522732896
transform 1 0 4344 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_38
timestamp 1522732896
transform 1 0 4424 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_2_0
timestamp 1522732896
transform 1 0 4616 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1522732896
transform 1 0 4632 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_2
timestamp 1522732896
transform 1 0 4648 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_46
timestamp 1522732896
transform 1 0 4664 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_213
timestamp 1522732896
transform -1 0 4920 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_214
timestamp 1522732896
transform -1 0 4984 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_154
timestamp 1522732896
transform 1 0 4984 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_62
timestamp 1522732896
transform -1 0 5096 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_39
timestamp 1522732896
transform -1 0 5144 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_67
timestamp 1522732896
transform -1 0 5176 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_64
timestamp 1522732896
transform -1 0 5368 0 -1 1410
box 0 0 192 200
use BUFX4  BUFX4_73
timestamp 1522732896
transform 1 0 5368 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_233
timestamp 1522732896
transform 1 0 5432 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_234
timestamp 1522732896
transform -1 0 5560 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_157
timestamp 1522732896
transform -1 0 5608 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_54
timestamp 1522732896
transform -1 0 5800 0 -1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_59
timestamp 1522732896
transform -1 0 5992 0 -1 1410
box 0 0 192 200
use AOI22X1  AOI22X1_35
timestamp 1522732896
transform -1 0 6072 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_48
timestamp 1522732896
transform -1 0 6264 0 -1 1410
box 0 0 192 200
use FILL  FILL_7_1
timestamp 1522732896
transform -1 0 6280 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_2
timestamp 1522732896
transform -1 0 6296 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_2
timestamp 1522732896
transform 1 0 8 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_56
timestamp 1522732896
transform 1 0 72 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_15
timestamp 1522732896
transform 1 0 120 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_16
timestamp 1522732896
transform 1 0 168 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_67
timestamp 1522732896
transform -1 0 264 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_23
timestamp 1522732896
transform 1 0 264 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_48
timestamp 1522732896
transform 1 0 312 0 1 1010
box 0 0 48 200
use INVX1  INVX1_34
timestamp 1522732896
transform -1 0 392 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_70
timestamp 1522732896
transform -1 0 440 0 1 1010
box 0 0 48 200
use INVX2  INVX2_1
timestamp 1522732896
transform 1 0 440 0 1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_18
timestamp 1522732896
transform -1 0 536 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1522732896
transform -1 0 600 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_2
timestamp 1522732896
transform 1 0 600 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_2
timestamp 1522732896
transform -1 0 712 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_1
timestamp 1522732896
transform -1 0 776 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_84
timestamp 1522732896
transform 1 0 776 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_71
timestamp 1522732896
transform 1 0 840 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_57
timestamp 1522732896
transform -1 0 952 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_64
timestamp 1522732896
transform -1 0 1000 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_87
timestamp 1522732896
transform -1 0 1048 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_78
timestamp 1522732896
transform -1 0 1096 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_76
timestamp 1522732896
transform -1 0 1144 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_68
timestamp 1522732896
transform 1 0 1144 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_48
timestamp 1522732896
transform -1 0 1272 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_3
timestamp 1522732896
transform -1 0 1336 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_81
timestamp 1522732896
transform 1 0 1336 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_128
timestamp 1522732896
transform 1 0 1384 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_94
timestamp 1522732896
transform -1 0 1512 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_56
timestamp 1522732896
transform 1 0 1512 0 1 1010
box 0 0 48 200
use INVX2  INVX2_25
timestamp 1522732896
transform 1 0 1560 0 1 1010
box 0 0 32 200
use FILL  FILL_5_0_0
timestamp 1522732896
transform 1 0 1592 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1522732896
transform 1 0 1608 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_2
timestamp 1522732896
transform 1 0 1624 0 1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_42
timestamp 1522732896
transform 1 0 1640 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_54
timestamp 1522732896
transform -1 0 1752 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_103
timestamp 1522732896
transform 1 0 1752 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_206
timestamp 1522732896
transform 1 0 1800 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_47
timestamp 1522732896
transform 1 0 1848 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_62
timestamp 1522732896
transform 1 0 1896 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_75
timestamp 1522732896
transform -1 0 2008 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_14
timestamp 1522732896
transform 1 0 2008 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_207
timestamp 1522732896
transform -1 0 2120 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_54
timestamp 1522732896
transform -1 0 2168 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_60
timestamp 1522732896
transform -1 0 2216 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_40
timestamp 1522732896
transform -1 0 2264 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_20
timestamp 1522732896
transform 1 0 2264 0 1 1010
box 0 0 64 200
use INVX4  INVX4_3
timestamp 1522732896
transform -1 0 2376 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_62
timestamp 1522732896
transform -1 0 2440 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_74
timestamp 1522732896
transform -1 0 2504 0 1 1010
box 0 0 64 200
use OAI22X1  OAI22X1_8
timestamp 1522732896
transform 1 0 2504 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_80
timestamp 1522732896
transform -1 0 2632 0 1 1010
box 0 0 48 200
use INVX1  INVX1_74
timestamp 1522732896
transform 1 0 2632 0 1 1010
box 0 0 32 200
use AND2X2  AND2X2_35
timestamp 1522732896
transform 1 0 2664 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_5
timestamp 1522732896
transform -1 0 2792 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_71
timestamp 1522732896
transform -1 0 2840 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_82
timestamp 1522732896
transform 1 0 2840 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_13
timestamp 1522732896
transform -1 0 2952 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1522732896
transform 1 0 2952 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_97
timestamp 1522732896
transform -1 0 3064 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_166
timestamp 1522732896
transform 1 0 3064 0 1 1010
box 0 0 64 200
use FILL  FILL_5_1_0
timestamp 1522732896
transform -1 0 3144 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1522732896
transform -1 0 3160 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_2
timestamp 1522732896
transform -1 0 3176 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_36
timestamp 1522732896
transform -1 0 3368 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_152
timestamp 1522732896
transform 1 0 3368 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_200
timestamp 1522732896
transform -1 0 3480 0 1 1010
box 0 0 64 200
use INVX1  INVX1_41
timestamp 1522732896
transform -1 0 3512 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_69
timestamp 1522732896
transform -1 0 3560 0 1 1010
box 0 0 48 200
use INVX1  INVX1_120
timestamp 1522732896
transform 1 0 3560 0 1 1010
box 0 0 32 200
use INVX1  INVX1_110
timestamp 1522732896
transform 1 0 3592 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_61
timestamp 1522732896
transform -1 0 3816 0 1 1010
box 0 0 192 200
use OAI22X1  OAI22X1_40
timestamp 1522732896
transform 1 0 3816 0 1 1010
box 0 0 80 200
use INVX1  INVX1_130
timestamp 1522732896
transform 1 0 3896 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_66
timestamp 1522732896
transform 1 0 3928 0 1 1010
box 0 0 192 200
use INVX1  INVX1_68
timestamp 1522732896
transform 1 0 4120 0 1 1010
box 0 0 32 200
use AOI21X1  AOI21X1_80
timestamp 1522732896
transform 1 0 4152 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_60
timestamp 1522732896
transform 1 0 4216 0 1 1010
box 0 0 64 200
use INVX1  INVX1_131
timestamp 1522732896
transform -1 0 4312 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_85
timestamp 1522732896
transform 1 0 4312 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_159
timestamp 1522732896
transform 1 0 4360 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_55
timestamp 1522732896
transform 1 0 4408 0 1 1010
box 0 0 192 200
use OAI22X1  OAI22X1_38
timestamp 1522732896
transform 1 0 4600 0 1 1010
box 0 0 80 200
use FILL  FILL_5_2_0
timestamp 1522732896
transform -1 0 4696 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1522732896
transform -1 0 4712 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_2
timestamp 1522732896
transform -1 0 4728 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_258
timestamp 1522732896
transform -1 0 4792 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_257
timestamp 1522732896
transform -1 0 4856 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_39
timestamp 1522732896
transform 1 0 4856 0 1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_250
timestamp 1522732896
transform -1 0 5000 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_181
timestamp 1522732896
transform 1 0 5000 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_260
timestamp 1522732896
transform -1 0 5112 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_136
timestamp 1522732896
transform -1 0 5176 0 1 1010
box 0 0 64 200
use INVX1  INVX1_142
timestamp 1522732896
transform -1 0 5208 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_177
timestamp 1522732896
transform -1 0 5256 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_161
timestamp 1522732896
transform 1 0 5256 0 1 1010
box 0 0 48 200
use INVX1  INVX1_140
timestamp 1522732896
transform -1 0 5336 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_155
timestamp 1522732896
transform -1 0 5384 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_158
timestamp 1522732896
transform 1 0 5384 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_160
timestamp 1522732896
transform 1 0 5432 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_162
timestamp 1522732896
transform 1 0 5480 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_38
timestamp 1522732896
transform 1 0 5528 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_161
timestamp 1522732896
transform 1 0 5608 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_159
timestamp 1522732896
transform -1 0 5704 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_244
timestamp 1522732896
transform 1 0 5704 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_220
timestamp 1522732896
transform 1 0 5768 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_219
timestamp 1522732896
transform -1 0 5896 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_168
timestamp 1522732896
transform -1 0 5944 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_162
timestamp 1522732896
transform 1 0 5944 0 1 1010
box 0 0 48 200
use INVX1  INVX1_137
timestamp 1522732896
transform 1 0 5992 0 1 1010
box 0 0 32 200
use AOI22X1  AOI22X1_36
timestamp 1522732896
transform -1 0 6104 0 1 1010
box 0 0 80 200
use INVX1  INVX1_106
timestamp 1522732896
transform -1 0 6136 0 1 1010
box 0 0 32 200
use OR2X2  OR2X2_19
timestamp 1522732896
transform -1 0 6200 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_419
timestamp 1522732896
transform 1 0 6200 0 1 1010
box 0 0 64 200
use FILL  FILL_6_1
timestamp 1522732896
transform 1 0 6264 0 1 1010
box 0 0 16 200
use FILL  FILL_6_2
timestamp 1522732896
transform 1 0 6280 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_1
timestamp 1522732896
transform 1 0 8 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_15
timestamp 1522732896
transform 1 0 56 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_75
timestamp 1522732896
transform 1 0 104 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_11
timestamp 1522732896
transform -1 0 200 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_12
timestamp 1522732896
transform -1 0 248 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_9
timestamp 1522732896
transform -1 0 296 0 -1 1010
box 0 0 48 200
use AND2X2  AND2X2_1
timestamp 1522732896
transform 1 0 296 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_59
timestamp 1522732896
transform 1 0 360 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_2
timestamp 1522732896
transform 1 0 408 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_13
timestamp 1522732896
transform -1 0 488 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_1
timestamp 1522732896
transform -1 0 536 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_61
timestamp 1522732896
transform -1 0 584 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_51
timestamp 1522732896
transform -1 0 648 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_94
timestamp 1522732896
transform -1 0 696 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_19
timestamp 1522732896
transform 1 0 696 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_21
timestamp 1522732896
transform 1 0 760 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_18
timestamp 1522732896
transform -1 0 872 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_77
timestamp 1522732896
transform 1 0 872 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_211
timestamp 1522732896
transform -1 0 968 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_91
timestamp 1522732896
transform 1 0 968 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_101
timestamp 1522732896
transform 1 0 1032 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_47
timestamp 1522732896
transform -1 0 1112 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_3
timestamp 1522732896
transform 1 0 1112 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_39
timestamp 1522732896
transform -1 0 1208 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_40
timestamp 1522732896
transform -1 0 1240 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_54
timestamp 1522732896
transform -1 0 1304 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_5
timestamp 1522732896
transform -1 0 1352 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_99
timestamp 1522732896
transform 1 0 1352 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_51
timestamp 1522732896
transform 1 0 1416 0 -1 1010
box 0 0 32 200
use INVX2  INVX2_27
timestamp 1522732896
transform 1 0 1448 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_93
timestamp 1522732896
transform -1 0 1544 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_45
timestamp 1522732896
transform 1 0 1544 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_0_0
timestamp 1522732896
transform 1 0 1608 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1522732896
transform 1 0 1624 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_2
timestamp 1522732896
transform 1 0 1640 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_60
timestamp 1522732896
transform 1 0 1656 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_142
timestamp 1522732896
transform -1 0 1784 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_69
timestamp 1522732896
transform -1 0 1848 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_89
timestamp 1522732896
transform -1 0 1912 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_67
timestamp 1522732896
transform 1 0 1912 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_50
timestamp 1522732896
transform 1 0 1976 0 -1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_95
timestamp 1522732896
transform -1 0 2056 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_78
timestamp 1522732896
transform 1 0 2056 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_88
timestamp 1522732896
transform 1 0 2104 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_95
timestamp 1522732896
transform 1 0 2152 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_94
timestamp 1522732896
transform 1 0 2216 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_120
timestamp 1522732896
transform -1 0 2344 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_108
timestamp 1522732896
transform -1 0 2392 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_14
timestamp 1522732896
transform 1 0 2392 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_36
timestamp 1522732896
transform 1 0 2456 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_70
timestamp 1522732896
transform 1 0 2488 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_68
timestamp 1522732896
transform -1 0 2600 0 -1 1010
box 0 0 48 200
use OR2X2  OR2X2_6
timestamp 1522732896
transform 1 0 2600 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_47
timestamp 1522732896
transform -1 0 2728 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_72
timestamp 1522732896
transform -1 0 2776 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_1
timestamp 1522732896
transform -1 0 2840 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_53
timestamp 1522732896
transform 1 0 2840 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_113
timestamp 1522732896
transform 1 0 2872 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_114
timestamp 1522732896
transform -1 0 3000 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_50
timestamp 1522732896
transform 1 0 3000 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_49
timestamp 1522732896
transform 1 0 3064 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_1_0
timestamp 1522732896
transform -1 0 3144 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1522732896
transform -1 0 3160 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_2
timestamp 1522732896
transform -1 0 3176 0 -1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_52
timestamp 1522732896
transform -1 0 3240 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_14
timestamp 1522732896
transform 1 0 3240 0 -1 1010
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_67
timestamp 1522732896
transform 1 0 3320 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_265
timestamp 1522732896
transform -1 0 3576 0 -1 1010
box 0 0 64 200
use INVX2  INVX2_30
timestamp 1522732896
transform 1 0 3576 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_60
timestamp 1522732896
transform -1 0 3800 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_245
timestamp 1522732896
transform 1 0 3800 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_46
timestamp 1522732896
transform -1 0 3912 0 -1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_62
timestamp 1522732896
transform -1 0 4104 0 -1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_47
timestamp 1522732896
transform 1 0 4104 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_7
timestamp 1522732896
transform 1 0 4152 0 -1 1010
box 0 0 48 200
use AND2X2  AND2X2_9
timestamp 1522732896
transform -1 0 4264 0 -1 1010
box 0 0 64 200
use BUFX2  BUFX2_9
timestamp 1522732896
transform 1 0 4264 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_8
timestamp 1522732896
transform 1 0 4312 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_105
timestamp 1522732896
transform -1 0 4424 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_16
timestamp 1522732896
transform 1 0 4424 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_70
timestamp 1522732896
transform -1 0 4536 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_72
timestamp 1522732896
transform -1 0 4600 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_15
timestamp 1522732896
transform 1 0 4600 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_2_0
timestamp 1522732896
transform 1 0 4664 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1522732896
transform 1 0 4680 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_2
timestamp 1522732896
transform 1 0 4696 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_229
timestamp 1522732896
transform 1 0 4712 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_90
timestamp 1522732896
transform -1 0 4824 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_79
timestamp 1522732896
transform 1 0 4824 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_180
timestamp 1522732896
transform 1 0 4888 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_254
timestamp 1522732896
transform -1 0 5000 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_252
timestamp 1522732896
transform -1 0 5064 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_177
timestamp 1522732896
transform -1 0 5112 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_178
timestamp 1522732896
transform 1 0 5112 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_247
timestamp 1522732896
transform 1 0 5160 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_249
timestamp 1522732896
transform 1 0 5224 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_248
timestamp 1522732896
transform -1 0 5352 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_203
timestamp 1522732896
transform -1 0 5416 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_134
timestamp 1522732896
transform -1 0 5448 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_255
timestamp 1522732896
transform 1 0 5448 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_165
timestamp 1522732896
transform 1 0 5512 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_256
timestamp 1522732896
transform -1 0 5624 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_175
timestamp 1522732896
transform -1 0 5672 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_30
timestamp 1522732896
transform -1 0 5736 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_78
timestamp 1522732896
transform -1 0 5800 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_28
timestamp 1522732896
transform 1 0 5800 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_138
timestamp 1522732896
transform 1 0 5864 0 -1 1010
box 0 0 32 200
use INVX1  INVX1_136
timestamp 1522732896
transform 1 0 5896 0 -1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_171
timestamp 1522732896
transform -1 0 5976 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_222
timestamp 1522732896
transform 1 0 5976 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_51
timestamp 1522732896
transform -1 0 6232 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_442
timestamp 1522732896
transform 1 0 6232 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_8
timestamp 1522732896
transform 1 0 8 0 1 610
box 0 0 48 200
use INVX1  INVX1_5
timestamp 1522732896
transform 1 0 56 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_5
timestamp 1522732896
transform -1 0 136 0 1 610
box 0 0 48 200
use INVX1  INVX1_7
timestamp 1522732896
transform 1 0 136 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_10
timestamp 1522732896
transform -1 0 216 0 1 610
box 0 0 48 200
use INVX1  INVX1_6
timestamp 1522732896
transform 1 0 216 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_6
timestamp 1522732896
transform -1 0 296 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_22
timestamp 1522732896
transform 1 0 296 0 1 610
box 0 0 48 200
use INVX1  INVX1_4
timestamp 1522732896
transform 1 0 344 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_4
timestamp 1522732896
transform -1 0 424 0 1 610
box 0 0 48 200
use OR2X2  OR2X2_1
timestamp 1522732896
transform 1 0 424 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_9
timestamp 1522732896
transform -1 0 536 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_59
timestamp 1522732896
transform -1 0 584 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_4
timestamp 1522732896
transform 1 0 584 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_50
timestamp 1522732896
transform 1 0 632 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_52
timestamp 1522732896
transform -1 0 728 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_16
timestamp 1522732896
transform 1 0 728 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_67
timestamp 1522732896
transform 1 0 776 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_157
timestamp 1522732896
transform 1 0 824 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_51
timestamp 1522732896
transform 1 0 888 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_156
timestamp 1522732896
transform -1 0 1000 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_308
timestamp 1522732896
transform -1 0 1064 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_44
timestamp 1522732896
transform -1 0 1128 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_48
timestamp 1522732896
transform 1 0 1128 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_52
timestamp 1522732896
transform 1 0 1176 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_23
timestamp 1522732896
transform -1 0 1288 0 1 610
box 0 0 48 200
use INVX2  INVX2_10
timestamp 1522732896
transform 1 0 1288 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_112
timestamp 1522732896
transform 1 0 1320 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_53
timestamp 1522732896
transform 1 0 1368 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_74
timestamp 1522732896
transform -1 0 1464 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_48
timestamp 1522732896
transform 1 0 1464 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_49
timestamp 1522732896
transform 1 0 1528 0 1 610
box 0 0 48 200
use FILL  FILL_3_0_0
timestamp 1522732896
transform -1 0 1592 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1522732896
transform -1 0 1608 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_2
timestamp 1522732896
transform -1 0 1624 0 1 610
box 0 0 16 200
use INVX1  INVX1_35
timestamp 1522732896
transform -1 0 1656 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_55
timestamp 1522732896
transform 1 0 1656 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_54
timestamp 1522732896
transform -1 0 1784 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_96
timestamp 1522732896
transform -1 0 1848 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_51
timestamp 1522732896
transform 1 0 1848 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_51
timestamp 1522732896
transform 1 0 1912 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_82
timestamp 1522732896
transform 1 0 1976 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_83
timestamp 1522732896
transform -1 0 2104 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1522732896
transform 1 0 2104 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_112
timestamp 1522732896
transform 1 0 2168 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_121
timestamp 1522732896
transform 1 0 2216 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_122
timestamp 1522732896
transform 1 0 2280 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_88
timestamp 1522732896
transform 1 0 2344 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_57
timestamp 1522732896
transform 1 0 2408 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1522732896
transform -1 0 2536 0 1 610
box 0 0 64 200
use NOR3X1  NOR3X1_6
timestamp 1522732896
transform 1 0 2536 0 1 610
box 0 0 128 200
use NOR2X1  NOR2X1_127
timestamp 1522732896
transform 1 0 2664 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_119
timestamp 1522732896
transform -1 0 2776 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_109
timestamp 1522732896
transform -1 0 2824 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_57
timestamp 1522732896
transform -1 0 2872 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_98
timestamp 1522732896
transform 1 0 2872 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_68
timestamp 1522732896
transform 1 0 2936 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_8
timestamp 1522732896
transform 1 0 3000 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_88
timestamp 1522732896
transform -1 0 3128 0 1 610
box 0 0 64 200
use FILL  FILL_3_1_0
timestamp 1522732896
transform 1 0 3128 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1522732896
transform 1 0 3144 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_2
timestamp 1522732896
transform 1 0 3160 0 1 610
box 0 0 16 200
use BUFX2  BUFX2_41
timestamp 1522732896
transform 1 0 3176 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_89
timestamp 1522732896
transform 1 0 3224 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_111
timestamp 1522732896
transform 1 0 3272 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_25
timestamp 1522732896
transform 1 0 3320 0 1 610
box 0 0 80 200
use AOI22X1  AOI22X1_16
timestamp 1522732896
transform 1 0 3400 0 1 610
box 0 0 80 200
use INVX1  INVX1_45
timestamp 1522732896
transform 1 0 3480 0 1 610
box 0 0 32 200
use AOI22X1  AOI22X1_17
timestamp 1522732896
transform 1 0 3512 0 1 610
box 0 0 80 200
use OAI21X1  OAI21X1_124
timestamp 1522732896
transform 1 0 3592 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_8
timestamp 1522732896
transform 1 0 3656 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_15
timestamp 1522732896
transform 1 0 3720 0 1 610
box 0 0 80 200
use BUFX4  BUFX4_67
timestamp 1522732896
transform -1 0 3864 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_99
timestamp 1522732896
transform 1 0 3864 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_101
timestamp 1522732896
transform -1 0 3976 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_98
timestamp 1522732896
transform 1 0 3976 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_143
timestamp 1522732896
transform 1 0 4024 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_142
timestamp 1522732896
transform -1 0 4152 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_58
timestamp 1522732896
transform 1 0 4152 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_55
timestamp 1522732896
transform 1 0 4200 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_47
timestamp 1522732896
transform 1 0 4248 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_10
timestamp 1522732896
transform -1 0 4376 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_56
timestamp 1522732896
transform 1 0 4376 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_41
timestamp 1522732896
transform 1 0 4440 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_89
timestamp 1522732896
transform -1 0 4536 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_37
timestamp 1522732896
transform 1 0 4536 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_97
timestamp 1522732896
transform 1 0 4600 0 1 610
box 0 0 48 200
use FILL  FILL_3_2_0
timestamp 1522732896
transform -1 0 4664 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1522732896
transform -1 0 4680 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_2
timestamp 1522732896
transform -1 0 4696 0 1 610
box 0 0 16 200
use INVX1  INVX1_44
timestamp 1522732896
transform -1 0 4728 0 1 610
box 0 0 32 200
use NAND3X1  NAND3X1_141
timestamp 1522732896
transform 1 0 4728 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_176
timestamp 1522732896
transform 1 0 4792 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_174
timestamp 1522732896
transform -1 0 4888 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_164
timestamp 1522732896
transform -1 0 4936 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_253
timestamp 1522732896
transform -1 0 5000 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_83
timestamp 1522732896
transform 1 0 5000 0 1 610
box 0 0 48 200
use INVX2  INVX2_29
timestamp 1522732896
transform 1 0 5048 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_107
timestamp 1522732896
transform -1 0 5128 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_34
timestamp 1522732896
transform -1 0 5208 0 1 610
box 0 0 80 200
use INVX1  INVX1_143
timestamp 1522732896
transform 1 0 5208 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_96
timestamp 1522732896
transform -1 0 5288 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_165
timestamp 1522732896
transform 1 0 5288 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_166
timestamp 1522732896
transform 1 0 5336 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_144
timestamp 1522732896
transform 1 0 5384 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_137
timestamp 1522732896
transform 1 0 5448 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_160
timestamp 1522732896
transform 1 0 5512 0 1 610
box 0 0 48 200
use OAI22X1  OAI22X1_37
timestamp 1522732896
transform -1 0 5640 0 1 610
box 0 0 80 200
use AOI21X1  AOI21X1_75
timestamp 1522732896
transform 1 0 5640 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_167
timestamp 1522732896
transform 1 0 5704 0 1 610
box 0 0 48 200
use INVX1  INVX1_135
timestamp 1522732896
transform 1 0 5752 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_246
timestamp 1522732896
transform -1 0 5848 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_139
timestamp 1522732896
transform -1 0 5912 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_98
timestamp 1522732896
transform 1 0 5912 0 1 610
box 0 0 48 200
use OR2X2  OR2X2_9
timestamp 1522732896
transform -1 0 6024 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_45
timestamp 1522732896
transform -1 0 6072 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_170
timestamp 1522732896
transform 1 0 6072 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_169
timestamp 1522732896
transform 1 0 6120 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_216
timestamp 1522732896
transform -1 0 6232 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_42
timestamp 1522732896
transform 1 0 6232 0 1 610
box 0 0 64 200
use DFFSR  DFFSR_6
timestamp 1522732896
transform 1 0 8 0 -1 610
box 0 0 352 200
use NOR2X1  NOR2X1_49
timestamp 1522732896
transform 1 0 360 0 -1 610
box 0 0 48 200
use INVX1  INVX1_3
timestamp 1522732896
transform 1 0 408 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_2
timestamp 1522732896
transform -1 0 488 0 -1 610
box 0 0 48 200
use INVX8  INVX8_1
timestamp 1522732896
transform -1 0 568 0 -1 610
box 0 0 80 200
use BUFX4  BUFX4_7
timestamp 1522732896
transform -1 0 632 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_50
timestamp 1522732896
transform -1 0 696 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_3
timestamp 1522732896
transform -1 0 744 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_59
timestamp 1522732896
transform 1 0 744 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_60
timestamp 1522732896
transform 1 0 808 0 -1 610
box 0 0 48 200
use MUX2X1  MUX2X1_7
timestamp 1522732896
transform -1 0 952 0 -1 610
box 0 0 96 200
use BUFX4  BUFX4_52
timestamp 1522732896
transform 1 0 952 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_13
timestamp 1522732896
transform 1 0 1016 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_1
timestamp 1522732896
transform 1 0 1080 0 -1 610
box 0 0 80 200
use NOR2X1  NOR2X1_63
timestamp 1522732896
transform -1 0 1208 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_63
timestamp 1522732896
transform 1 0 1208 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_62
timestamp 1522732896
transform -1 0 1336 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_78
timestamp 1522732896
transform -1 0 1400 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_108
timestamp 1522732896
transform 1 0 1400 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_5
timestamp 1522732896
transform 1 0 1464 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_50
timestamp 1522732896
transform 1 0 1528 0 -1 610
box 0 0 48 200
use FILL  FILL_2_0_0
timestamp 1522732896
transform 1 0 1576 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1522732896
transform 1 0 1592 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_2
timestamp 1522732896
transform 1 0 1608 0 -1 610
box 0 0 16 200
use INVX1  INVX1_37
timestamp 1522732896
transform 1 0 1624 0 -1 610
box 0 0 32 200
use OR2X2  OR2X2_3
timestamp 1522732896
transform 1 0 1656 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_125
timestamp 1522732896
transform -1 0 1768 0 -1 610
box 0 0 48 200
use MUX2X1  MUX2X1_8
timestamp 1522732896
transform -1 0 1864 0 -1 610
box 0 0 96 200
use NOR2X1  NOR2X1_122
timestamp 1522732896
transform 1 0 1864 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_76
timestamp 1522732896
transform -1 0 1976 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_81
timestamp 1522732896
transform 1 0 1976 0 -1 610
box 0 0 64 200
use INVX1  INVX1_56
timestamp 1522732896
transform -1 0 2072 0 -1 610
box 0 0 32 200
use INVX1  INVX1_57
timestamp 1522732896
transform -1 0 2104 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_106
timestamp 1522732896
transform 1 0 2104 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_107
timestamp 1522732896
transform -1 0 2232 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_76
timestamp 1522732896
transform -1 0 2280 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_77
timestamp 1522732896
transform -1 0 2344 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_77
timestamp 1522732896
transform -1 0 2392 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_104
timestamp 1522732896
transform 1 0 2392 0 -1 610
box 0 0 48 200
use AOI21X1  AOI21X1_43
timestamp 1522732896
transform -1 0 2504 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_81
timestamp 1522732896
transform 1 0 2504 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_80
timestamp 1522732896
transform -1 0 2632 0 -1 610
box 0 0 64 200
use INVX1  INVX1_59
timestamp 1522732896
transform -1 0 2664 0 -1 610
box 0 0 32 200
use BUFX4  BUFX4_12
timestamp 1522732896
transform 1 0 2664 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_117
timestamp 1522732896
transform 1 0 2728 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_53
timestamp 1522732896
transform -1 0 2856 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_75
timestamp 1522732896
transform 1 0 2856 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_88
timestamp 1522732896
transform -1 0 2952 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_87
timestamp 1522732896
transform 1 0 2952 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_86
timestamp 1522732896
transform 1 0 3016 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_86
timestamp 1522732896
transform -1 0 3128 0 -1 610
box 0 0 48 200
use FILL  FILL_2_1_0
timestamp 1522732896
transform 1 0 3128 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1522732896
transform 1 0 3144 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_2
timestamp 1522732896
transform 1 0 3160 0 -1 610
box 0 0 16 200
use AND2X2  AND2X2_24
timestamp 1522732896
transform 1 0 3176 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_87
timestamp 1522732896
transform 1 0 3240 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_128
timestamp 1522732896
transform -1 0 3352 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_63
timestamp 1522732896
transform 1 0 3352 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_89
timestamp 1522732896
transform -1 0 3480 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_72
timestamp 1522732896
transform 1 0 3480 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_94
timestamp 1522732896
transform 1 0 3544 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_113
timestamp 1522732896
transform 1 0 3592 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_120
timestamp 1522732896
transform 1 0 3640 0 -1 610
box 0 0 48 200
use OAI22X1  OAI22X1_6
timestamp 1522732896
transform 1 0 3688 0 -1 610
box 0 0 80 200
use OAI21X1  OAI21X1_127
timestamp 1522732896
transform 1 0 3768 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_7
timestamp 1522732896
transform 1 0 3832 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_65
timestamp 1522732896
transform 1 0 3896 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_44
timestamp 1522732896
transform -1 0 4024 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_108
timestamp 1522732896
transform 1 0 4024 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_59
timestamp 1522732896
transform -1 0 4136 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_93
timestamp 1522732896
transform -1 0 4184 0 -1 610
box 0 0 48 200
use MUX2X1  MUX2X1_21
timestamp 1522732896
transform 1 0 4184 0 -1 610
box 0 0 96 200
use AND2X2  AND2X2_19
timestamp 1522732896
transform -1 0 4344 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_27
timestamp 1522732896
transform -1 0 4408 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_58
timestamp 1522732896
transform -1 0 4472 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_70
timestamp 1522732896
transform -1 0 4536 0 -1 610
box 0 0 64 200
use NOR3X1  NOR3X1_5
timestamp 1522732896
transform 1 0 4536 0 -1 610
box 0 0 128 200
use FILL  FILL_2_2_0
timestamp 1522732896
transform 1 0 4664 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1522732896
transform 1 0 4680 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_2
timestamp 1522732896
transform 1 0 4696 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_83
timestamp 1522732896
transform 1 0 4712 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_43
timestamp 1522732896
transform 1 0 4760 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_112
timestamp 1522732896
transform -1 0 4888 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_86
timestamp 1522732896
transform 1 0 4888 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_29
timestamp 1522732896
transform -1 0 5000 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_59
timestamp 1522732896
transform 1 0 5000 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_91
timestamp 1522732896
transform -1 0 5112 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_61
timestamp 1522732896
transform 1 0 5112 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_179
timestamp 1522732896
transform 1 0 5176 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_41
timestamp 1522732896
transform -1 0 5272 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_43
timestamp 1522732896
transform -1 0 5320 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_73
timestamp 1522732896
transform -1 0 5368 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_264
timestamp 1522732896
transform -1 0 5432 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_20
timestamp 1522732896
transform -1 0 5496 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_261
timestamp 1522732896
transform -1 0 5560 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_145
timestamp 1522732896
transform 1 0 5560 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_163
timestamp 1522732896
transform -1 0 5672 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_232
timestamp 1522732896
transform 1 0 5672 0 -1 610
box 0 0 64 200
use OAI22X1  OAI22X1_41
timestamp 1522732896
transform -1 0 5816 0 -1 610
box 0 0 80 200
use NOR2X1  NOR2X1_104
timestamp 1522732896
transform 1 0 5816 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_172
timestamp 1522732896
transform -1 0 5912 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_88
timestamp 1522732896
transform -1 0 5976 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_175
timestamp 1522732896
transform 1 0 5976 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_221
timestamp 1522732896
transform 1 0 6024 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_76
timestamp 1522732896
transform 1 0 6088 0 -1 610
box 0 0 64 200
use INVX8  INVX8_6
timestamp 1522732896
transform 1 0 6152 0 -1 610
box 0 0 80 200
use BUFX4  BUFX4_40
timestamp 1522732896
transform -1 0 6296 0 -1 610
box 0 0 64 200
use DFFSR  DFFSR_2
timestamp 1522732896
transform -1 0 360 0 1 210
box 0 0 352 200
use DFFSR  DFFSR_1
timestamp 1522732896
transform -1 0 712 0 1 210
box 0 0 352 200
use DFFSR  DFFSR_5
timestamp 1522732896
transform -1 0 1064 0 1 210
box 0 0 352 200
use NAND2X1  NAND2X1_93
timestamp 1522732896
transform 1 0 1064 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_89
timestamp 1522732896
transform -1 0 1176 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_53
timestamp 1522732896
transform 1 0 1176 0 1 210
box 0 0 48 200
use INVX1  INVX1_54
timestamp 1522732896
transform 1 0 1224 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_49
timestamp 1522732896
transform 1 0 1256 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_79
timestamp 1522732896
transform 1 0 1320 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_11
timestamp 1522732896
transform 1 0 1384 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_50
timestamp 1522732896
transform 1 0 1448 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_110
timestamp 1522732896
transform 1 0 1512 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1522732896
transform 1 0 1576 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1522732896
transform 1 0 1592 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_2
timestamp 1522732896
transform 1 0 1608 0 1 210
box 0 0 16 200
use OAI21X1  OAI21X1_111
timestamp 1522732896
transform 1 0 1624 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_124
timestamp 1522732896
transform -1 0 1736 0 1 210
box 0 0 48 200
use AND2X2  AND2X2_25
timestamp 1522732896
transform 1 0 1736 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_85
timestamp 1522732896
transform -1 0 1864 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_109
timestamp 1522732896
transform -1 0 1928 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_45
timestamp 1522732896
transform 1 0 1928 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_52
timestamp 1522732896
transform 1 0 1992 0 1 210
box 0 0 48 200
use OR2X2  OR2X2_11
timestamp 1522732896
transform 1 0 2040 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_116
timestamp 1522732896
transform -1 0 2152 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_106
timestamp 1522732896
transform -1 0 2200 0 1 210
box 0 0 48 200
use AND2X2  AND2X2_23
timestamp 1522732896
transform -1 0 2264 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_12
timestamp 1522732896
transform 1 0 2264 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_69
timestamp 1522732896
transform 1 0 2328 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_61
timestamp 1522732896
transform -1 0 2440 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_116
timestamp 1522732896
transform 1 0 2440 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1522732896
transform 1 0 2504 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_126
timestamp 1522732896
transform -1 0 2600 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_86
timestamp 1522732896
transform 1 0 2600 0 1 210
box 0 0 64 200
use AOI21X1  AOI21X1_49
timestamp 1522732896
transform -1 0 2728 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_109
timestamp 1522732896
transform 1 0 2728 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_74
timestamp 1522732896
transform -1 0 2840 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_110
timestamp 1522732896
transform -1 0 2888 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_55
timestamp 1522732896
transform 1 0 2888 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_57
timestamp 1522732896
transform -1 0 3000 0 1 210
box 0 0 64 200
use AOI21X1  AOI21X1_48
timestamp 1522732896
transform 1 0 3000 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_113
timestamp 1522732896
transform -1 0 3112 0 1 210
box 0 0 48 200
use FILL  FILL_1_1_0
timestamp 1522732896
transform 1 0 3112 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1522732896
transform 1 0 3128 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_2
timestamp 1522732896
transform 1 0 3144 0 1 210
box 0 0 16 200
use NOR3X1  NOR3X1_9
timestamp 1522732896
transform 1 0 3160 0 1 210
box 0 0 128 200
use NOR3X1  NOR3X1_7
timestamp 1522732896
transform 1 0 3288 0 1 210
box 0 0 128 200
use OAI21X1  OAI21X1_115
timestamp 1522732896
transform 1 0 3416 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_119
timestamp 1522732896
transform -1 0 3528 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_84
timestamp 1522732896
transform 1 0 3528 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_121
timestamp 1522732896
transform 1 0 3592 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_61
timestamp 1522732896
transform 1 0 3640 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_125
timestamp 1522732896
transform -1 0 3768 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_83
timestamp 1522732896
transform -1 0 3832 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_123
timestamp 1522732896
transform -1 0 3896 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_60
timestamp 1522732896
transform 1 0 3896 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_24
timestamp 1522732896
transform 1 0 3960 0 1 210
box 0 0 80 200
use OAI22X1  OAI22X1_9
timestamp 1522732896
transform -1 0 4120 0 1 210
box 0 0 80 200
use NOR3X1  NOR3X1_11
timestamp 1522732896
transform 1 0 4120 0 1 210
box 0 0 128 200
use OAI22X1  OAI22X1_10
timestamp 1522732896
transform 1 0 4248 0 1 210
box 0 0 80 200
use NAND2X1  NAND2X1_115
timestamp 1522732896
transform 1 0 4328 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_114
timestamp 1522732896
transform 1 0 4376 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_120
timestamp 1522732896
transform -1 0 4472 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_64
timestamp 1522732896
transform 1 0 4472 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_76
timestamp 1522732896
transform 1 0 4536 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_19
timestamp 1522732896
transform -1 0 4680 0 1 210
box 0 0 80 200
use FILL  FILL_1_2_0
timestamp 1522732896
transform 1 0 4680 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1522732896
transform 1 0 4696 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_2
timestamp 1522732896
transform 1 0 4712 0 1 210
box 0 0 16 200
use NAND3X1  NAND3X1_71
timestamp 1522732896
transform 1 0 4728 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_23
timestamp 1522732896
transform -1 0 4872 0 1 210
box 0 0 80 200
use NOR2X1  NOR2X1_106
timestamp 1522732896
transform 1 0 4872 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_73
timestamp 1522732896
transform -1 0 4968 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_71
timestamp 1522732896
transform 1 0 4968 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_72
timestamp 1522732896
transform 1 0 5016 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_92
timestamp 1522732896
transform -1 0 5112 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_85
timestamp 1522732896
transform -1 0 5160 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_97
timestamp 1522732896
transform -1 0 5224 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_82
timestamp 1522732896
transform 1 0 5224 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_65
timestamp 1522732896
transform -1 0 5320 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_138
timestamp 1522732896
transform 1 0 5320 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_20
timestamp 1522732896
transform -1 0 5464 0 1 210
box 0 0 80 200
use NAND3X1  NAND3X1_69
timestamp 1522732896
transform 1 0 5464 0 1 210
box 0 0 64 200
use AOI21X1  AOI21X1_46
timestamp 1522732896
transform -1 0 5592 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_262
timestamp 1522732896
transform 1 0 5592 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_21
timestamp 1522732896
transform 1 0 5656 0 1 210
box 0 0 80 200
use NOR2X1  NOR2X1_184
timestamp 1522732896
transform -1 0 5784 0 1 210
box 0 0 48 200
use AOI21X1  AOI21X1_77
timestamp 1522732896
transform 1 0 5784 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_182
timestamp 1522732896
transform -1 0 5896 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_102
timestamp 1522732896
transform 1 0 5896 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_173
timestamp 1522732896
transform -1 0 5992 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_103
timestamp 1522732896
transform -1 0 6056 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_215
timestamp 1522732896
transform -1 0 6120 0 1 210
box 0 0 64 200
use INVX1  INVX1_133
timestamp 1522732896
transform 1 0 6120 0 1 210
box 0 0 32 200
use NAND3X1  NAND3X1_140
timestamp 1522732896
transform 1 0 6152 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_42
timestamp 1522732896
transform -1 0 6264 0 1 210
box 0 0 48 200
use FILL  FILL_2_1
timestamp 1522732896
transform 1 0 6264 0 1 210
box 0 0 16 200
use FILL  FILL_2_2
timestamp 1522732896
transform 1 0 6280 0 1 210
box 0 0 16 200
use DFFSR  DFFSR_4
timestamp 1522732896
transform 1 0 8 0 -1 210
box 0 0 352 200
use DFFSR  DFFSR_3
timestamp 1522732896
transform -1 0 712 0 -1 210
box 0 0 352 200
use INVX8  INVX8_5
timestamp 1522732896
transform -1 0 792 0 -1 210
box 0 0 80 200
use BUFX4  BUFX4_74
timestamp 1522732896
transform 1 0 792 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_52
timestamp 1522732896
transform 1 0 856 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_90
timestamp 1522732896
transform 1 0 920 0 -1 210
box 0 0 64 200
use INVX1  INVX1_38
timestamp 1522732896
transform 1 0 984 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_53
timestamp 1522732896
transform -1 0 1080 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_62
timestamp 1522732896
transform 1 0 1080 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_65
timestamp 1522732896
transform 1 0 1128 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_61
timestamp 1522732896
transform -1 0 1240 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_68
timestamp 1522732896
transform 1 0 1240 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_117
timestamp 1522732896
transform 1 0 1288 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_73
timestamp 1522732896
transform -1 0 1400 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_115
timestamp 1522732896
transform -1 0 1448 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_118
timestamp 1522732896
transform -1 0 1496 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_12
timestamp 1522732896
transform 1 0 1496 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_64
timestamp 1522732896
transform 1 0 1560 0 -1 210
box 0 0 48 200
use FILL  FILL_0_0_0
timestamp 1522732896
transform -1 0 1624 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1522732896
transform -1 0 1640 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_2
timestamp 1522732896
transform -1 0 1656 0 -1 210
box 0 0 16 200
use OR2X2  OR2X2_4
timestamp 1522732896
transform -1 0 1720 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_123
timestamp 1522732896
transform 1 0 1720 0 -1 210
box 0 0 48 200
use INVX1  INVX1_58
timestamp 1522732896
transform -1 0 1800 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_117
timestamp 1522732896
transform -1 0 1848 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_79
timestamp 1522732896
transform 1 0 1848 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_82
timestamp 1522732896
transform -1 0 1976 0 -1 210
box 0 0 64 200
use INVX1  INVX1_52
timestamp 1522732896
transform 1 0 1976 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_107
timestamp 1522732896
transform -1 0 2056 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_55
timestamp 1522732896
transform 1 0 2056 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_58
timestamp 1522732896
transform 1 0 2120 0 -1 210
box 0 0 64 200
use INVX1  INVX1_42
timestamp 1522732896
transform -1 0 2216 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_79
timestamp 1522732896
transform 1 0 2216 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_81
timestamp 1522732896
transform -1 0 2312 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_69
timestamp 1522732896
transform 1 0 2312 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_66
timestamp 1522732896
transform 1 0 2360 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_80
timestamp 1522732896
transform 1 0 2424 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_56
timestamp 1522732896
transform 1 0 2472 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_75
timestamp 1522732896
transform 1 0 2536 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_111
timestamp 1522732896
transform -1 0 2648 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_110
timestamp 1522732896
transform -1 0 2696 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_21
timestamp 1522732896
transform -1 0 2760 0 -1 210
box 0 0 64 200
use INVX1  INVX1_49
timestamp 1522732896
transform -1 0 2792 0 -1 210
box 0 0 32 200
use NAND3X1  NAND3X1_78
timestamp 1522732896
transform 1 0 2792 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_126
timestamp 1522732896
transform 1 0 2856 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_10
timestamp 1522732896
transform -1 0 2984 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_77
timestamp 1522732896
transform -1 0 3048 0 -1 210
box 0 0 64 200
use INVX1  INVX1_55
timestamp 1522732896
transform 1 0 3048 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_114
timestamp 1522732896
transform -1 0 3128 0 -1 210
box 0 0 48 200
use FILL  FILL_0_1_0
timestamp 1522732896
transform -1 0 3144 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1522732896
transform -1 0 3160 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_2
timestamp 1522732896
transform -1 0 3176 0 -1 210
box 0 0 16 200
use NOR3X1  NOR3X1_10
timestamp 1522732896
transform -1 0 3304 0 -1 210
box 0 0 128 200
use AND2X2  AND2X2_22
timestamp 1522732896
transform 1 0 3304 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_80
timestamp 1522732896
transform 1 0 3368 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_118
timestamp 1522732896
transform 1 0 3432 0 -1 210
box 0 0 48 200
use AOI21X1  AOI21X1_39
timestamp 1522732896
transform -1 0 3544 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_41
timestamp 1522732896
transform -1 0 3608 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_17
timestamp 1522732896
transform -1 0 3672 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_95
timestamp 1522732896
transform 1 0 3672 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_18
timestamp 1522732896
transform -1 0 3784 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_116
timestamp 1522732896
transform -1 0 3832 0 -1 210
box 0 0 48 200
use AOI22X1  AOI22X1_18
timestamp 1522732896
transform 1 0 3832 0 -1 210
box 0 0 80 200
use NAND2X1  NAND2X1_119
timestamp 1522732896
transform 1 0 3912 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_101
timestamp 1522732896
transform 1 0 3960 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_68
timestamp 1522732896
transform -1 0 4072 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_102
timestamp 1522732896
transform -1 0 4136 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_100
timestamp 1522732896
transform 1 0 4136 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_91
timestamp 1522732896
transform 1 0 4184 0 -1 210
box 0 0 48 200
use AOI21X1  AOI21X1_47
timestamp 1522732896
transform 1 0 4232 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_22
timestamp 1522732896
transform 1 0 4296 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_67
timestamp 1522732896
transform -1 0 4440 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_90
timestamp 1522732896
transform -1 0 4488 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_84
timestamp 1522732896
transform -1 0 4536 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_105
timestamp 1522732896
transform 1 0 4536 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_87
timestamp 1522732896
transform -1 0 4632 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_105
timestamp 1522732896
transform -1 0 4680 0 -1 210
box 0 0 48 200
use FILL  FILL_0_2_0
timestamp 1522732896
transform -1 0 4696 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1522732896
transform -1 0 4712 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_2
timestamp 1522732896
transform -1 0 4728 0 -1 210
box 0 0 16 200
use NOR3X1  NOR3X1_8
timestamp 1522732896
transform -1 0 4856 0 -1 210
box 0 0 128 200
use NOR2X1  NOR2X1_66
timestamp 1522732896
transform -1 0 4904 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_66
timestamp 1522732896
transform -1 0 4968 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_65
timestamp 1522732896
transform 1 0 4968 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_43
timestamp 1522732896
transform 1 0 5032 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_263
timestamp 1522732896
transform 1 0 5080 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_183
timestamp 1522732896
transform 1 0 5144 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_103
timestamp 1522732896
transform 1 0 5192 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_44
timestamp 1522732896
transform -1 0 5288 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_104
timestamp 1522732896
transform -1 0 5352 0 -1 210
box 0 0 64 200
use INVX1  INVX1_149
timestamp 1522732896
transform -1 0 5384 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_227
timestamp 1522732896
transform 1 0 5384 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_41
timestamp 1522732896
transform 1 0 5448 0 -1 210
box 0 0 64 200
use INVX1  INVX1_109
timestamp 1522732896
transform 1 0 5512 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_49
timestamp 1522732896
transform -1 0 5736 0 -1 210
box 0 0 192 200
use INVX1  INVX1_205
timestamp 1522732896
transform -1 0 5768 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_53
timestamp 1522732896
transform -1 0 5960 0 -1 210
box 0 0 192 200
use MUX2X1  MUX2X1_35
timestamp 1522732896
transform 1 0 5960 0 -1 210
box 0 0 96 200
use BUFX4  BUFX4_37
timestamp 1522732896
transform 1 0 6056 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_129
timestamp 1522732896
transform 1 0 6120 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_242
timestamp 1522732896
transform -1 0 6232 0 -1 210
box 0 0 48 200
use INVX1  INVX1_191
timestamp 1522732896
transform -1 0 6264 0 -1 210
box 0 0 32 200
use FILL  FILL_1_1
timestamp 1522732896
transform -1 0 6280 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1522732896
transform -1 0 6296 0 -1 210
box 0 0 16 200
<< labels >>
flabel metal4 1576 -40 1624 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 3112 -40 3160 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 400 4640 400 4640 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal3 -16 1520 -16 1520 7 FreeSans 24 0 0 0 reset
port 3 nsew
flabel metal2 640 4640 640 4640 3 FreeSans 24 90 0 0 DI<0>
port 4 nsew
flabel metal3 -16 1320 -16 1320 7 FreeSans 24 0 0 0 DI<1>
port 5 nsew
flabel metal2 2752 4640 2752 4640 3 FreeSans 24 90 0 0 DI<2>
port 6 nsew
flabel metal3 -16 4520 -16 4520 7 FreeSans 24 0 0 0 DI<3>
port 7 nsew
flabel space 3200 4640 3200 4640 3 FreeSans 24 90 0 0 DI<4>
port 8 nsew
flabel metal2 1056 4640 1056 4640 3 FreeSans 24 90 0 0 DI<5>
port 9 nsew
flabel space 3200 -20 3200 -20 7 FreeSans 24 270 0 0 DI<6>
port 10 nsew
flabel space 3280 -20 3280 -20 7 FreeSans 24 270 0 0 DI<7>
port 11 nsew
flabel metal2 2864 4640 2864 4640 3 FreeSans 24 90 0 0 IRQ
port 12 nsew
flabel metal2 2464 4640 2464 4640 3 FreeSans 24 90 0 0 NMI
port 13 nsew
flabel metal3 -16 2300 -16 2300 7 FreeSans 24 0 0 0 RDY
port 14 nsew
flabel metal2 592 4640 592 4640 3 FreeSans 24 90 0 0 AB<0>
port 15 nsew
flabel metal2 1840 4640 1840 4640 3 FreeSans 24 90 0 0 AB<1>
port 16 nsew
flabel metal2 1904 4640 1904 4640 3 FreeSans 24 90 0 0 AB<2>
port 17 nsew
flabel metal2 2096 4640 2096 4640 3 FreeSans 24 90 0 0 AB<3>
port 18 nsew
flabel metal2 1168 4640 1168 4640 3 FreeSans 24 90 0 0 AB<4>
port 19 nsew
flabel metal2 1760 4640 1760 4640 3 FreeSans 24 90 0 0 AB<5>
port 20 nsew
flabel metal2 2000 4640 2000 4640 3 FreeSans 24 90 0 0 AB<6>
port 21 nsew
flabel metal2 880 4640 880 4640 3 FreeSans 24 90 0 0 AB<7>
port 22 nsew
flabel metal2 2240 4640 2240 4640 3 FreeSans 24 90 0 0 AB<8>
port 23 nsew
flabel metal2 752 4640 752 4640 3 FreeSans 24 90 0 0 AB<9>
port 24 nsew
flabel metal2 1408 4640 1408 4640 3 FreeSans 24 90 0 0 AB<10>
port 25 nsew
flabel metal2 2160 4640 2160 4640 3 FreeSans 24 90 0 0 AB<11>
port 26 nsew
flabel metal2 1712 4640 1712 4640 3 FreeSans 24 90 0 0 AB<12>
port 27 nsew
flabel metal2 1952 4640 1952 4640 3 FreeSans 24 90 0 0 AB<13>
port 28 nsew
flabel metal2 1632 4640 1632 4640 3 FreeSans 24 90 0 0 AB<14>
port 29 nsew
flabel metal2 2032 4640 2032 4640 3 FreeSans 24 90 0 0 AB<15>
port 30 nsew
flabel metal2 2512 4640 2512 4640 3 FreeSans 24 90 0 0 DO<0>
port 31 nsew
flabel metal2 3504 4640 3504 4640 3 FreeSans 24 90 0 0 DO<1>
port 32 nsew
flabel metal2 2640 4640 2640 4640 3 FreeSans 24 90 0 0 DO<2>
port 33 nsew
flabel metal2 3120 4640 3120 4640 3 FreeSans 24 90 0 0 DO<3>
port 34 nsew
flabel metal2 3248 4640 3248 4640 3 FreeSans 24 90 0 0 DO<4>
port 35 nsew
flabel metal2 3312 4640 3312 4640 3 FreeSans 24 90 0 0 DO<5>
port 36 nsew
flabel metal2 2912 4640 2912 4640 3 FreeSans 24 90 0 0 DO<6>
port 37 nsew
flabel metal2 2800 4640 2800 4640 3 FreeSans 24 90 0 0 DO<7>
port 38 nsew
flabel metal2 3248 -20 3248 -20 7 FreeSans 24 270 0 0 WE
port 39 nsew
<< end >>
